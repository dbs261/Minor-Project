`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.04.2022 22:35:14
// Design Name: 
// Module Name: Multiplier
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Multiplier(
    input [31:0] X,
    input [31:0] Y,
    output [63:0] Z
    );
wire X0Y0, X0Y1, X0Y2, X0Y3, X0Y4, X0Y5, X0Y6, X0Y7, X0Y8, X0Y9, X0Y10, X0Y11, X0Y12, X0Y13, X0Y14, X0Y15, X0Y16, X0Y17, X0Y18, X0Y19, X0Y20, X0Y21, X0Y22, X0Y23, X0Y24, X0Y25, X0Y26, X0Y27, X0Y28, X0Y29, X0Y30, X0Y31;
wire X1Y0, X1Y1, X1Y2, X1Y3, X1Y4, X1Y5, X1Y6, X1Y7, X1Y8, X1Y9, X1Y10, X1Y11, X1Y12, X1Y13, X1Y14, X1Y15, X1Y16, X1Y17, X1Y18, X1Y19, X1Y20, X1Y21, X1Y22, X1Y23, X1Y24, X1Y25, X1Y26, X1Y27, X1Y28, X1Y29, X1Y30, X1Y31;
wire X2Y0, X2Y1, X2Y2, X2Y3, X2Y4, X2Y5, X2Y6, X2Y7, X2Y8, X2Y9, X2Y10, X2Y11, X2Y12, X2Y13, X2Y14, X2Y15, X2Y16, X2Y17, X2Y18, X2Y19, X2Y20, X2Y21, X2Y22, X2Y23, X2Y24, X2Y25, X2Y26, X2Y27, X2Y28, X2Y29, X2Y30, X2Y31;
    wire X3Y0, X3Y1, X3Y2, X3Y3, X3Y4, X3Y5, X3Y6, X3Y7, X3Y8, X3Y9, X3Y10, X3Y11, X3Y12, X3Y13, X3Y14, X3Y15, X3Y16, X3Y17, X3Y18, X3Y19, X3Y20, X3Y21, X3Y22, X3Y23, X3Y24, X3Y25, X3Y26, X3Y27, X3Y28, X3Y29, X3Y30, X3Y31;
    wire X4Y0, X4Y1, X4Y2, X4Y3, X4Y4, X4Y5, X4Y6, X4Y7, X4Y8, X4Y9, X4Y10, X4Y11, X4Y12, X4Y13, X4Y14, X4Y15, X4Y16, X4Y17, X4Y18, X4Y19, X4Y20, X4Y21, X4Y22, X4Y23, X4Y24, X4Y25, X4Y26, X4Y27, X4Y28, X4Y29, X4Y30, X4Y31;
    wire X5Y0, X5Y1, X5Y2, X5Y3, X5Y4, X5Y5, X5Y6, X5Y7, X5Y8, X5Y9, X5Y10, X5Y11, X5Y12, X5Y13, X5Y14, X5Y15, X5Y16, X5Y17, X5Y18, X5Y19, X5Y20, X5Y21, X5Y22, X5Y23, X5Y24, X5Y25, X5Y26, X5Y27, X5Y28, X5Y29, X5Y30, X5Y31;
    wire X6Y0, X6Y1, X6Y2, X6Y3, X6Y4, X6Y5, X6Y6, X6Y7, X6Y8, X6Y9, X6Y10, X6Y11, X6Y12, X6Y13, X6Y14, X6Y15, X6Y16, X6Y17, X6Y18, X6Y19, X6Y20, X6Y21, X6Y22, X6Y23, X6Y24, X6Y25, X6Y26, X6Y27, X6Y28, X6Y29, X6Y30, X6Y31;
    wire X7Y0, X7Y1, X7Y2, X7Y3, X7Y4, X7Y5, X7Y6, X7Y7, X7Y8, X7Y9, X7Y10, X7Y11, X7Y12, X7Y13, X7Y14, X7Y15, X7Y16, X7Y17, X7Y18, X7Y19, X7Y20, X7Y21, X7Y22, X7Y23, X7Y24, X7Y25, X7Y26, X7Y27, X7Y28, X7Y29, X7Y30, X7Y31;
    wire X8Y0, X8Y1, X8Y2, X8Y3, X8Y4, X8Y5, X8Y6, X8Y7, X8Y8, X8Y9, X8Y10, X8Y11, X8Y12, X8Y13, X8Y14, X8Y15, X8Y16, X8Y17, X8Y18, X8Y19, X8Y20, X8Y21, X8Y22, X8Y23, X8Y24, X8Y25, X8Y26, X8Y27, X8Y28, X8Y29, X8Y30, X8Y31;
    wire X9Y0, X9Y1, X9Y2, X9Y3, X9Y4, X9Y5, X9Y6, X9Y7, X9Y8, X9Y9, X9Y10, X9Y11, X9Y12, X9Y13, X9Y14, X9Y15, X9Y16, X9Y17, X9Y18, X9Y19, X9Y20, X9Y21, X9Y22, X9Y23, X9Y24, X9Y25, X9Y26, X9Y27, X9Y28, X9Y29, X9Y30, X9Y31;
    wire X10Y0, X10Y1, X10Y2, X10Y3, X10Y4, X10Y5, X10Y6, X10Y7, X10Y8, X10Y9, X10Y10, X10Y11, X10Y12, X10Y13, X10Y14, X10Y15, X10Y16, X10Y17, X10Y18, X10Y19, X10Y20, X10Y21, X10Y22, X10Y23, X10Y24, X10Y25, X10Y26, X10Y27, X10Y28, X10Y29, X10Y30, X10Y31;
    wire X11Y0, X11Y1, X11Y2, X11Y3, X11Y4, X11Y5, X11Y6, X11Y7, X11Y8, X11Y9, X11Y10, X11Y11, X11Y12, X11Y13, X11Y14, X11Y15, X11Y16, X11Y17, X11Y18, X11Y19, X11Y20, X11Y21, X11Y22, X11Y23, X11Y24, X11Y25, X11Y26, X11Y27, X11Y28, X11Y29, X11Y30, X11Y31;
    wire X12Y0, X12Y1, X12Y2, X12Y3, X12Y4, X12Y5, X12Y6, X12Y7, X12Y8, X12Y9, X12Y10, X12Y11, X12Y12, X12Y13, X12Y14, X12Y15, X12Y16, X12Y17, X12Y18, X12Y19, X12Y20, X12Y21, X12Y22, X12Y23, X12Y24, X12Y25, X12Y26, X12Y27, X12Y28, X12Y29, X12Y30, X12Y31;
    wire X13Y0, X13Y1, X13Y2, X13Y3, X13Y4, X13Y5, X13Y6, X13Y7, X13Y8, X13Y9, X13Y10, X13Y11, X13Y12, X13Y13, X13Y14, X13Y15, X13Y16, X13Y17, X13Y18, X13Y19, X13Y20, X13Y21, X13Y22, X13Y23, X13Y24, X13Y25, X13Y26, X13Y27, X13Y28, X13Y29, X13Y30, X13Y31;
    wire X14Y0, X14Y1, X14Y2, X14Y3, X14Y4, X14Y5, X14Y6, X14Y7, X14Y8, X14Y9, X14Y10, X14Y11, X14Y12, X14Y13, X14Y14, X14Y15, X14Y16, X14Y17, X14Y18, X14Y19, X14Y20, X14Y21, X14Y22, X14Y23, X14Y24, X14Y25, X14Y26, X14Y27, X14Y28, X14Y29, X14Y30, X14Y31;
    wire X15Y0, X15Y1, X15Y2, X15Y3, X15Y4, X15Y5, X15Y6, X15Y7, X15Y8, X15Y9, X15Y10, X15Y11, X15Y12, X15Y13, X15Y14, X15Y15, X15Y16, X15Y17, X15Y18, X15Y19, X15Y20, X15Y21, X15Y22, X15Y23, X15Y24, X15Y25, X15Y26, X15Y27, X15Y28, X15Y29, X15Y30, X15Y31;
    wire X16Y0, X16Y1, X16Y2, X16Y3, X16Y4, X16Y5, X16Y6, X16Y7, X16Y8, X16Y9, X16Y10, X16Y11, X16Y12, X16Y13, X16Y14, X16Y15, X16Y16, X16Y17, X16Y18, X16Y19, X16Y20, X16Y21, X16Y22, X16Y23, X16Y24, X16Y25, X16Y26, X16Y27, X16Y28, X16Y29, X16Y30, X16Y31;
    wire X17Y0, X17Y1, X17Y2, X17Y3, X17Y4, X17Y5, X17Y6, X17Y7, X17Y8, X17Y9, X17Y10, X17Y11, X17Y12, X17Y13, X17Y14, X17Y15, X17Y16, X17Y17, X17Y18, X17Y19, X17Y20, X17Y21, X17Y22, X17Y23, X17Y24, X17Y25, X17Y26, X17Y27, X17Y28, X17Y29, X17Y30, X17Y31;
    wire X18Y0, X18Y1, X18Y2, X18Y3, X18Y4, X18Y5, X18Y6, X18Y7, X18Y8, X18Y9, X18Y10, X18Y11, X18Y12, X18Y13, X18Y14, X18Y15, X18Y16, X18Y17, X18Y18, X18Y19, X18Y20, X18Y21, X18Y22, X18Y23, X18Y24, X18Y25, X18Y26, X18Y27, X18Y28, X18Y29, X18Y30, X18Y31;
    wire X19Y0, X19Y1, X19Y2, X19Y3, X19Y4, X19Y5, X19Y6, X19Y7, X19Y8, X19Y9, X19Y10, X19Y11, X19Y12, X19Y13, X19Y14, X19Y15, X19Y16, X19Y17, X19Y18, X19Y19, X19Y20, X19Y21, X19Y22, X19Y23, X19Y24, X19Y25, X19Y26, X19Y27, X19Y28, X19Y29, X19Y30, X19Y31;
    wire X20Y0, X20Y1, X20Y2, X20Y3, X20Y4, X20Y5, X20Y6, X20Y7, X20Y8, X20Y9, X20Y10, X20Y11, X20Y12, X20Y13, X20Y14, X20Y15, X20Y16, X20Y17, X20Y18, X20Y19, X20Y20, X20Y21, X20Y22, X20Y23, X20Y24, X20Y25, X20Y26, X20Y27, X20Y28, X20Y29, X20Y30, X20Y31;
    wire X21Y0, X21Y1, X21Y2, X21Y3, X21Y4, X21Y5, X21Y6, X21Y7, X21Y8, X21Y9, X21Y10, X21Y11, X21Y12, X21Y13, X21Y14, X21Y15, X21Y16, X21Y17, X21Y18, X21Y19, X21Y20, X21Y21, X21Y22, X21Y23, X21Y24, X21Y25, X21Y26, X21Y27, X21Y28, X21Y29, X21Y30, X21Y31;
    wire X22Y0, X22Y1, X22Y2, X22Y3, X22Y4, X22Y5, X22Y6, X22Y7, X22Y8, X22Y9, X22Y10, X22Y11, X22Y12, X22Y13, X22Y14, X22Y15, X22Y16, X22Y17, X22Y18, X22Y19, X22Y20, X22Y21, X22Y22, X22Y23, X22Y24, X22Y25, X22Y26, X22Y27, X22Y28, X22Y29, X22Y30, X22Y31;
    wire X23Y0, X23Y1, X23Y2, X23Y3, X23Y4, X23Y5, X23Y6, X23Y7, X23Y8, X23Y9, X23Y10, X23Y11, X23Y12, X23Y13, X23Y14, X23Y15, X23Y16, X23Y17, X23Y18, X23Y19, X23Y20, X23Y21, X23Y22, X23Y23, X23Y24, X23Y25, X23Y26, X23Y27, X23Y28, X23Y29, X23Y30, X23Y31;
    wire X24Y0, X24Y1, X24Y2, X24Y3, X24Y4, X24Y5, X24Y6, X24Y7, X24Y8, X24Y9, X24Y10, X24Y11, X24Y12, X24Y13, X24Y14, X24Y15, X24Y16, X24Y17, X24Y18, X24Y19, X24Y20, X24Y21, X24Y22, X24Y23, X24Y24, X24Y25, X24Y26, X24Y27, X24Y28, X24Y29, X24Y30, X24Y31;
    wire X25Y0, X25Y1, X25Y2, X25Y3, X25Y4, X25Y5, X25Y6, X25Y7, X25Y8, X25Y9, X25Y10, X25Y11, X25Y12, X25Y13, X25Y14, X25Y15, X25Y16, X25Y17, X25Y18, X25Y19, X25Y20, X25Y21, X25Y22, X25Y23, X25Y24, X25Y25, X25Y26, X25Y27, X25Y28, X25Y29, X25Y30, X25Y31;
    wire X26Y0, X26Y1, X26Y2, X26Y3, X26Y4, X26Y5, X26Y6, X26Y7, X26Y8, X26Y9, X26Y10, X26Y11, X26Y12, X26Y13, X26Y14, X26Y15, X26Y16, X26Y17, X26Y18, X26Y19, X26Y20, X26Y21, X26Y22, X26Y23, X26Y24, X26Y25, X26Y26, X26Y27, X26Y28, X26Y29, X26Y30, X26Y31;
    wire X27Y0, X27Y1, X27Y2, X27Y3, X27Y4, X27Y5, X27Y6, X27Y7, X27Y8, X27Y9, X27Y10, X27Y11, X27Y12, X27Y13, X27Y14, X27Y15, X27Y16, X27Y17, X27Y18, X27Y19, X27Y20, X27Y21, X27Y22, X27Y23, X27Y24, X27Y25, X27Y26, X27Y27, X27Y28, X27Y29, X27Y30, X27Y31;
    wire X28Y0, X28Y1, X28Y2, X28Y3, X28Y4, X28Y5, X28Y6, X28Y7, X28Y8, X28Y9, X28Y10, X28Y11, X28Y12, X28Y13, X28Y14, X28Y15, X28Y16, X28Y17, X28Y18, X28Y19, X28Y20, X28Y21, X28Y22, X28Y23, X28Y24, X28Y25, X28Y26, X28Y27, X28Y28, X28Y29, X28Y30, X28Y31;
    wire X29Y0, X29Y1, X29Y2, X29Y3, X29Y4, X29Y5, X29Y6, X29Y7, X29Y8, X29Y9, X29Y10, X29Y11, X29Y12, X29Y13, X29Y14, X29Y15, X29Y16, X29Y17, X29Y18, X29Y19, X29Y20, X29Y21, X29Y22, X29Y23, X29Y24, X29Y25, X29Y26, X29Y27, X29Y28, X29Y29, X29Y30, X29Y31;
    wire X30Y0, X30Y1, X30Y2, X30Y3, X30Y4, X30Y5, X30Y6, X30Y7, X30Y8, X30Y9, X30Y10, X30Y11, X30Y12, X30Y13, X30Y14, X30Y15, X30Y16, X30Y17, X30Y18, X30Y19, X30Y20, X30Y21, X30Y22, X30Y23, X30Y24, X30Y25, X30Y26, X30Y27, X30Y28, X30Y29, X30Y30, X30Y31;
    wire X31Y0, X31Y1, X31Y2, X31Y3, X31Y4, X31Y5, X31Y6, X31Y7, X31Y8, X31Y9, X31Y10, X31Y11, X31Y12, X31Y13, X31Y14, X31Y15, X31Y16, X31Y17, X31Y18, X31Y19, X31Y20, X31Y21, X31Y22, X31Y23, X31Y24, X31Y25, X31Y26, X31Y27, X31Y28, X31Y29, X31Y30, X31Y31;

wire c1_0, c1_1, c1_2, c1_3, c1_4, c1_5, c1_6, c1_7, c1_8, c1_9, c1_10, c1_11, c1_12, c1_13, c1_14, c1_15, c1_16, c1_17, c1_18, c1_19, c1_20, c1_21, c1_22, c1_23, c1_24, c1_25, c1_26, c1_27, c1_28, c1_29, c1_30, c1_31;
wire c2_0, c2_1, c2_2, c2_3, c2_4, c2_5, c2_6, c2_7, c2_8, c2_9, c2_10, c2_11, c2_12, c2_13, c2_14, c2_15, c2_16, c2_17, c2_18, c2_19, c2_20, c2_21, c2_22, c2_23, c2_24, c2_25, c2_26, c2_27, c2_28, c2_29, c2_30, c2_31;
wire c3_0, c3_1, c3_2, c3_3, c3_4, c3_5, c3_6, c3_7, c3_8, c3_9, c3_10, c3_11, c3_12, c3_13, c3_14, c3_15, c3_16, c3_17, c3_18, c3_19, c3_20, c3_21, c3_22, c3_23, c3_24, c3_25, c3_26, c3_27, c3_28, c3_29, c3_30, c3_31;
wire c4_0, c4_1, c4_2, c4_3, c4_4, c4_5, c4_6, c4_7, c4_8, c4_9, c4_10, c4_11, c4_12, c4_13, c4_14, c4_15, c4_16, c4_17, c4_18, c4_19, c4_20, c4_21, c4_22, c4_23, c4_24, c4_25, c4_26, c4_27, c4_28, c4_29, c4_30, c4_31;
wire c5_0, c5_1, c5_2, c5_3, c5_4, c5_5, c5_6, c5_7, c5_8, c5_9, c5_10, c5_11, c5_12, c5_13, c5_14, c5_15, c5_16, c5_17, c5_18, c5_19, c5_20, c5_21, c5_22, c5_23, c5_24, c5_25, c5_26, c5_27, c5_28, c5_29, c5_30, c5_31;
wire c6_0, c6_1, c6_2, c6_3, c6_4, c6_5, c6_6, c6_7, c6_8, c6_9, c6_10, c6_11, c6_12, c6_13, c6_14, c6_15, c6_16, c6_17, c6_18, c6_19, c6_20, c6_21, c6_22, c6_23, c6_24, c6_25, c6_26, c6_27, c6_28, c6_29, c6_30, c6_31;
wire c7_0, c7_1, c7_2, c7_3, c7_4, c7_5, c7_6, c7_7, c7_8, c7_9, c7_10, c7_11, c7_12, c7_13, c7_14, c7_15, c7_16, c7_17, c7_18, c7_19, c7_20, c7_21, c7_22, c7_23, c7_24, c7_25, c7_26, c7_27, c7_28, c7_29, c7_30, c7_31;
wire c8_0, c8_1, c8_2, c8_3, c8_4, c8_5, c8_6, c8_7, c8_8, c8_9, c8_10, c8_11, c8_12, c8_13, c8_14, c8_15, c8_16, c8_17, c8_18, c8_19, c8_20, c8_21, c8_22, c8_23, c8_24, c8_25, c8_26, c8_27, c8_28, c8_29, c8_30, c8_31;
wire c9_0, c9_1, c9_2, c9_3, c9_4, c9_5, c9_6, c9_7, c9_8, c9_9, c9_10, c9_11, c9_12, c9_13, c9_14, c9_15, c9_16, c9_17, c9_18, c9_19, c9_20, c9_21, c9_22, c9_23, c9_24, c9_25, c9_26, c9_27, c9_28, c9_29, c9_30, c9_31;
wire c10_0, c10_1, c10_2, c10_3, c10_4, c10_5, c10_6, c10_7, c10_8, c10_9, c10_10, c10_11, c10_12, c10_13, c10_14, c10_15, c10_16, c10_17, c10_18, c10_19, c10_20, c10_21, c10_22, c10_23, c10_24, c10_25, c10_26, c10_27, c10_28, c10_29, c10_30, c10_31;
wire c11_0, c11_1, c11_2, c11_3, c11_4, c11_5, c11_6, c11_7, c11_8, c11_9, c11_10, c11_11, c11_12, c11_13, c11_14, c11_15, c11_16, c11_17, c11_18, c11_19, c11_20, c11_21, c11_22, c11_23, c11_24, c11_25, c11_26, c11_27, c11_28, c11_29, c11_30, c11_31;
wire c12_0, c12_1, c12_2, c12_3, c12_4, c12_5, c12_6, c12_7, c12_8, c12_9, c12_10, c12_11, c12_12, c12_13, c12_14, c12_15, c12_16, c12_17, c12_18, c12_19, c12_20, c12_21, c12_22, c12_23, c12_24, c12_25, c12_26, c12_27, c12_28, c12_29, c12_30, c12_31;
wire c13_0, c13_1, c13_2, c13_3, c13_4, c13_5, c13_6, c13_7, c13_8, c13_9, c13_10, c13_11, c13_12, c13_13, c13_14, c13_15, c13_16, c13_17, c13_18, c13_19, c13_20, c13_21, c13_22, c13_23, c13_24, c13_25, c13_26, c13_27, c13_28, c13_29, c13_30, c13_31;
wire c14_0, c14_1, c14_2, c14_3, c14_4, c14_5, c14_6, c14_7, c14_8, c14_9, c14_10, c14_11, c14_12, c14_13, c14_14, c14_15, c14_16, c14_17, c14_18, c14_19, c14_20, c14_21, c14_22, c14_23, c14_24, c14_25, c14_26, c14_27, c14_28, c14_29, c14_30, c14_31;
wire c15_0, c15_1, c15_2, c15_3, c15_4, c15_5, c15_6, c15_7, c15_8, c15_9, c15_10, c15_11, c15_12, c15_13, c15_14, c15_15, c15_16, c15_17, c15_18, c15_19, c15_20, c15_21, c15_22, c15_23, c15_24, c15_25, c15_26, c15_27, c15_28, c15_29, c15_30, c15_31;
wire c16_0, c16_1, c16_2, c16_3, c16_4, c16_5, c16_6, c16_7, c16_8, c16_9, c16_10, c16_11, c16_12, c16_13, c16_14, c16_15, c16_16, c16_17, c16_18, c16_19, c16_20, c16_21, c16_22, c16_23, c16_24, c16_25, c16_26, c16_27, c16_28, c16_29, c16_30, c16_31;
wire c17_0, c17_1, c17_2, c17_3, c17_4, c17_5, c17_6, c17_7, c17_8, c17_9, c17_10, c17_11, c17_12, c17_13, c17_14, c17_15, c17_16, c17_17, c17_18, c17_19, c17_20, c17_21, c17_22, c17_23, c17_24, c17_25, c17_26, c17_27, c17_28, c17_29, c17_30, c17_31;
wire c18_0, c18_1, c18_2, c18_3, c18_4, c18_5, c18_6, c18_7, c18_8, c18_9, c18_10, c18_11, c18_12, c18_13, c18_14, c18_15, c18_16, c18_17, c18_18, c18_19, c18_20, c18_21, c18_22, c18_23, c18_24, c18_25, c18_26, c18_27, c18_28, c18_29, c18_30, c18_31;
wire c19_0, c19_1, c19_2, c19_3, c19_4, c19_5, c19_6, c19_7, c19_8, c19_9, c19_10, c19_11, c19_12, c19_13, c19_14, c19_15, c19_16, c19_17, c19_18, c19_19, c19_20, c19_21, c19_22, c19_23, c19_24, c19_25, c19_26, c19_27, c19_28, c19_29, c19_30, c19_31;
wire c20_0, c20_1, c20_2, c20_3, c20_4, c20_5, c20_6, c20_7, c20_8, c20_9, c20_10, c20_11, c20_12, c20_13, c20_14, c20_15, c20_16, c20_17, c20_18, c20_19, c20_20, c20_21, c20_22, c20_23, c20_24, c20_25, c20_26, c20_27, c20_28, c20_29, c20_30, c20_31;
wire c21_0, c21_1, c21_2, c21_3, c21_4, c21_5, c21_6, c21_7, c21_8, c21_9, c21_10, c21_11, c21_12, c21_13, c21_14, c21_15, c21_16, c21_17, c21_18, c21_19, c21_20, c21_21, c21_22, c21_23, c21_24, c21_25, c21_26, c21_27, c21_28, c21_29, c21_30, c21_31;
wire c22_0, c22_1, c22_2, c22_3, c22_4, c22_5, c22_6, c22_7, c22_8, c22_9, c22_10, c22_11, c22_12, c22_13, c22_14, c22_15, c22_16, c22_17, c22_18, c22_19, c22_20, c22_21, c22_22, c22_23, c22_24, c22_25, c22_26, c22_27, c22_28, c22_29, c22_30, c22_31;
wire c23_0, c23_1, c23_2, c23_3, c23_4, c23_5, c23_6, c23_7, c23_8, c23_9, c23_10, c23_11, c23_12, c23_13, c23_14, c23_15, c23_16, c23_17, c23_18, c23_19, c23_20, c23_21, c23_22, c23_23, c23_24, c23_25, c23_26, c23_27, c23_28, c23_29, c23_30, c23_31;
wire c24_0, c24_1, c24_2, c24_3, c24_4, c24_5, c24_6, c24_7, c24_8, c24_9, c24_10, c24_11, c24_12, c24_13, c24_14, c24_15, c24_16, c24_17, c24_18, c24_19, c24_20, c24_21, c24_22, c24_23, c24_24, c24_25, c24_26, c24_27, c24_28, c24_29, c24_30, c24_31;
wire c25_0, c25_1, c25_2, c25_3, c25_4, c25_5, c25_6, c25_7, c25_8, c25_9, c25_10, c25_11, c25_12, c25_13, c25_14, c25_15, c25_16, c25_17, c25_18, c25_19, c25_20, c25_21, c25_22, c25_23, c25_24, c25_25, c25_26, c25_27, c25_28, c25_29, c25_30, c25_31;
wire c26_0, c26_1, c26_2, c26_3, c26_4, c26_5, c26_6, c26_7, c26_8, c26_9, c26_10, c26_11, c26_12, c26_13, c26_14, c26_15, c26_16, c26_17, c26_18, c26_19, c26_20, c26_21, c26_22, c26_23, c26_24, c26_25, c26_26, c26_27, c26_28, c26_29, c26_30, c26_31;
wire c27_0, c27_1, c27_2, c27_3, c27_4, c27_5, c27_6, c27_7, c27_8, c27_9, c27_10, c27_11, c27_12, c27_13, c27_14, c27_15, c27_16, c27_17, c27_18, c27_19, c27_20, c27_21, c27_22, c27_23, c27_24, c27_25, c27_26, c27_27, c27_28, c27_29, c27_30, c27_31;
wire c28_0, c28_1, c28_2, c28_3, c28_4, c28_5, c28_6, c28_7, c28_8, c28_9, c28_10, c28_11, c28_12, c28_13, c28_14, c28_15, c28_16, c28_17, c28_18, c28_19, c28_20, c28_21, c28_22, c28_23, c28_24, c28_25, c28_26, c28_27, c28_28, c28_29, c28_30, c28_31;
wire c29_0, c29_1, c29_2, c29_3, c29_4, c29_5, c29_6, c29_7, c29_8, c29_9, c29_10, c29_11, c29_12, c29_13, c29_14, c29_15, c29_16, c29_17, c29_18, c29_19, c29_20, c29_21, c29_22, c29_23, c29_24, c29_25, c29_26, c29_27, c29_28, c29_29, c29_30, c29_31;
wire c30_0, c30_1, c30_2, c30_3, c30_4, c30_5, c30_6, c30_7, c30_8, c30_9, c30_10, c30_11, c30_12, c30_13, c30_14, c30_15, c30_16, c30_17, c30_18, c30_19, c30_20, c30_21, c30_22, c30_23, c30_24, c30_25, c30_26, c30_27, c30_28, c30_29, c30_30, c30_31;
wire c31_0, c31_1, c31_2, c31_3, c31_4, c31_5, c31_6, c31_7, c31_8, c31_9, c31_10, c31_11, c31_12, c31_13, c31_14, c31_15, c31_16, c31_17, c31_18, c31_19, c31_20, c31_21, c31_22, c31_23, c31_24, c31_25, c31_26, c31_27, c31_28, c31_29, c31_30, c31_31;
wire c0_31;

wire z1_0, z1_1, z1_2, z1_3, z1_4, z1_5, z1_6, z1_7, z1_8, z1_9, z1_10, z1_11, z1_12, z1_13, z1_14, z1_15, z1_16, z1_17, z1_18, z1_19, z1_20, z1_21, z1_22, z1_23, z1_24, z1_25, z1_26, z1_27, z1_28, z1_29, z1_30, z1_31;
wire z2_0, z2_1, z2_2, z2_3, z2_4, z2_5, z2_6, z2_7, z2_8, z2_9, z2_10, z2_11, z2_12, z2_13, z2_14, z2_15, z2_16, z2_17, z2_18, z2_19, z2_20, z2_21, z2_22, z2_23, z2_24, z2_25, z2_26, z2_27, z2_28, z2_29, z2_30, z2_31;
wire z3_0, z3_1, z3_2, z3_3, z3_4, z3_5, z3_6, z3_7, z3_8, z3_9, z3_10, z3_11, z3_12, z3_13, z3_14, z3_15, z3_16, z3_17, z3_18, z3_19, z3_20, z3_21, z3_22, z3_23, z3_24, z3_25, z3_26, z3_27, z3_28, z3_29, z3_30, z3_31;
wire z4_0, z4_1, z4_2, z4_3, z4_4, z4_5, z4_6, z4_7, z4_8, z4_9, z4_10, z4_11, z4_12, z4_13, z4_14, z4_15, z4_16, z4_17, z4_18, z4_19, z4_20, z4_21, z4_22, z4_23, z4_24, z4_25, z4_26, z4_27, z4_28, z4_29, z4_30, z4_31;
wire z5_0, z5_1, z5_2, z5_3, z5_4, z5_5, z5_6, z5_7, z5_8, z5_9, z5_10, z5_11, z5_12, z5_13, z5_14, z5_15, z5_16, z5_17, z5_18, z5_19, z5_20, z5_21, z5_22, z5_23, z5_24, z5_25, z5_26, z5_27, z5_28, z5_29, z5_30, z5_31;
wire z6_0, z6_1, z6_2, z6_3, z6_4, z6_5, z6_6, z6_7, z6_8, z6_9, z6_10, z6_11, z6_12, z6_13, z6_14, z6_15, z6_16, z6_17, z6_18, z6_19, z6_20, z6_21, z6_22, z6_23, z6_24, z6_25, z6_26, z6_27, z6_28, z6_29, z6_30, z6_31;
wire z7_0, z7_1, z7_2, z7_3, z7_4, z7_5, z7_6, z7_7, z7_8, z7_9, z7_10, z7_11, z7_12, z7_13, z7_14, z7_15, z7_16, z7_17, z7_18, z7_19, z7_20, z7_21, z7_22, z7_23, z7_24, z7_25, z7_26, z7_27, z7_28, z7_29, z7_30, z7_31;
wire z8_0, z8_1, z8_2, z8_3, z8_4, z8_5, z8_6, z8_7, z8_8, z8_9, z8_10, z8_11, z8_12, z8_13, z8_14, z8_15, z8_16, z8_17, z8_18, z8_19, z8_20, z8_21, z8_22, z8_23, z8_24, z8_25, z8_26, z8_27, z8_28, z8_29, z8_30, z8_31;
wire z9_0, z9_1, z9_2, z9_3, z9_4, z9_5, z9_6, z9_7, z9_8, z9_9, z9_10, z9_11, z9_12, z9_13, z9_14, z9_15, z9_16, z9_17, z9_18, z9_19, z9_20, z9_21, z9_22, z9_23, z9_24, z9_25, z9_26, z9_27, z9_28, z9_29, z9_30, z9_31;
wire z10_0, z10_1, z10_2, z10_3, z10_4, z10_5, z10_6, z10_7, z10_8, z10_9, z10_10, z10_11, z10_12, z10_13, z10_14, z10_15, z10_16, z10_17, z10_18, z10_19, z10_20, z10_21, z10_22, z10_23, z10_24, z10_25, z10_26, z10_27, z10_28, z10_29, z10_30, z10_31;
wire z11_0, z11_1, z11_2, z11_3, z11_4, z11_5, z11_6, z11_7, z11_8, z11_9, z11_10, z11_11, z11_12, z11_13, z11_14, z11_15, z11_16, z11_17, z11_18, z11_19, z11_20, z11_21, z11_22, z11_23, z11_24, z11_25, z11_26, z11_27, z11_28, z11_29, z11_30, z11_31;
wire z12_0, z12_1, z12_2, z12_3, z12_4, z12_5, z12_6, z12_7, z12_8, z12_9, z12_10, z12_11, z12_12, z12_13, z12_14, z12_15, z12_16, z12_17, z12_18, z12_19, z12_20, z12_21, z12_22, z12_23, z12_24, z12_25, z12_26, z12_27, z12_28, z12_29, z12_30, z12_31;
wire z13_0, z13_1, z13_2, z13_3, z13_4, z13_5, z13_6, z13_7, z13_8, z13_9, z13_10, z13_11, z13_12, z13_13, z13_14, z13_15, z13_16, z13_17, z13_18, z13_19, z13_20, z13_21, z13_22, z13_23, z13_24, z13_25, z13_26, z13_27, z13_28, z13_29, z13_30, z13_31;
wire z14_0, z14_1, z14_2, z14_3, z14_4, z14_5, z14_6, z14_7, z14_8, z14_9, z14_10, z14_11, z14_12, z14_13, z14_14, z14_15, z14_16, z14_17, z14_18, z14_19, z14_20, z14_21, z14_22, z14_23, z14_24, z14_25, z14_26, z14_27, z14_28, z14_29, z14_30, z14_31;
wire z15_0, z15_1, z15_2, z15_3, z15_4, z15_5, z15_6, z15_7, z15_8, z15_9, z15_10, z15_11, z15_12, z15_13, z15_14, z15_15, z15_16, z15_17, z15_18, z15_19, z15_20, z15_21, z15_22, z15_23, z15_24, z15_25, z15_26, z15_27, z15_28, z15_29, z15_30, z15_31;
wire z16_0, z16_1, z16_2, z16_3, z16_4, z16_5, z16_6, z16_7, z16_8, z16_9, z16_10, z16_11, z16_12, z16_13, z16_14, z16_15, z16_16, z16_17, z16_18, z16_19, z16_20, z16_21, z16_22, z16_23, z16_24, z16_25, z16_26, z16_27, z16_28, z16_29, z16_30, z16_31;
wire z17_0, z17_1, z17_2, z17_3, z17_4, z17_5, z17_6, z17_7, z17_8, z17_9, z17_10, z17_11, z17_12, z17_13, z17_14, z17_15, z17_16, z17_17, z17_18, z17_19, z17_20, z17_21, z17_22, z17_23, z17_24, z17_25, z17_26, z17_27, z17_28, z17_29, z17_30, z17_31;
wire z18_0, z18_1, z18_2, z18_3, z18_4, z18_5, z18_6, z18_7, z18_8, z18_9, z18_10, z18_11, z18_12, z18_13, z18_14, z18_15, z18_16, z18_17, z18_18, z18_19, z18_20, z18_21, z18_22, z18_23, z18_24, z18_25, z18_26, z18_27, z18_28, z18_29, z18_30, z18_31;
wire z19_0, z19_1, z19_2, z19_3, z19_4, z19_5, z19_6, z19_7, z19_8, z19_9, z19_10, z19_11, z19_12, z19_13, z19_14, z19_15, z19_16, z19_17, z19_18, z19_19, z19_20, z19_21, z19_22, z19_23, z19_24, z19_25, z19_26, z19_27, z19_28, z19_29, z19_30, z19_31;
wire z20_0, z20_1, z20_2, z20_3, z20_4, z20_5, z20_6, z20_7, z20_8, z20_9, z20_10, z20_11, z20_12, z20_13, z20_14, z20_15, z20_16, z20_17, z20_18, z20_19, z20_20, z20_21, z20_22, z20_23, z20_24, z20_25, z20_26, z20_27, z20_28, z20_29, z20_30, z20_31;
wire z21_0, z21_1, z21_2, z21_3, z21_4, z21_5, z21_6, z21_7, z21_8, z21_9, z21_10, z21_11, z21_12, z21_13, z21_14, z21_15, z21_16, z21_17, z21_18, z21_19, z21_20, z21_21, z21_22, z21_23, z21_24, z21_25, z21_26, z21_27, z21_28, z21_29, z21_30, z21_31;
wire z22_0, z22_1, z22_2, z22_3, z22_4, z22_5, z22_6, z22_7, z22_8, z22_9, z22_10, z22_11, z22_12, z22_13, z22_14, z22_15, z22_16, z22_17, z22_18, z22_19, z22_20, z22_21, z22_22, z22_23, z22_24, z22_25, z22_26, z22_27, z22_28, z22_29, z22_30, z22_31;
wire z23_0, z23_1, z23_2, z23_3, z23_4, z23_5, z23_6, z23_7, z23_8, z23_9, z23_10, z23_11, z23_12, z23_13, z23_14, z23_15, z23_16, z23_17, z23_18, z23_19, z23_20, z23_21, z23_22, z23_23, z23_24, z23_25, z23_26, z23_27, z23_28, z23_29, z23_30, z23_31;
wire z24_0, z24_1, z24_2, z24_3, z24_4, z24_5, z24_6, z24_7, z24_8, z24_9, z24_10, z24_11, z24_12, z24_13, z24_14, z24_15, z24_16, z24_17, z24_18, z24_19, z24_20, z24_21, z24_22, z24_23, z24_24, z24_25, z24_26, z24_27, z24_28, z24_29, z24_30, z24_31;
wire z25_0, z25_1, z25_2, z25_3, z25_4, z25_5, z25_6, z25_7, z25_8, z25_9, z25_10, z25_11, z25_12, z25_13, z25_14, z25_15, z25_16, z25_17, z25_18, z25_19, z25_20, z25_21, z25_22, z25_23, z25_24, z25_25, z25_26, z25_27, z25_28, z25_29, z25_30, z25_31;
wire z26_0, z26_1, z26_2, z26_3, z26_4, z26_5, z26_6, z26_7, z26_8, z26_9, z26_10, z26_11, z26_12, z26_13, z26_14, z26_15, z26_16, z26_17, z26_18, z26_19, z26_20, z26_21, z26_22, z26_23, z26_24, z26_25, z26_26, z26_27, z26_28, z26_29, z26_30, z26_31;
wire z27_0, z27_1, z27_2, z27_3, z27_4, z27_5, z27_6, z27_7, z27_8, z27_9, z27_10, z27_11, z27_12, z27_13, z27_14, z27_15, z27_16, z27_17, z27_18, z27_19, z27_20, z27_21, z27_22, z27_23, z27_24, z27_25, z27_26, z27_27, z27_28, z27_29, z27_30, z27_31;
wire z28_0, z28_1, z28_2, z28_3, z28_4, z28_5, z28_6, z28_7, z28_8, z28_9, z28_10, z28_11, z28_12, z28_13, z28_14, z28_15, z28_16, z28_17, z28_18, z28_19, z28_20, z28_21, z28_22, z28_23, z28_24, z28_25, z28_26, z28_27, z28_28, z28_29, z28_30, z28_31;
wire z29_0, z29_1, z29_2, z29_3, z29_4, z29_5, z29_6, z29_7, z29_8, z29_9, z29_10, z29_11, z29_12, z29_13, z29_14, z29_15, z29_16, z29_17, z29_18, z29_19, z29_20, z29_21, z29_22, z29_23, z29_24, z29_25, z29_26, z29_27, z29_28, z29_29, z29_30, z29_31;
wire z30_0, z30_1, z30_2, z30_3, z30_4, z30_5, z30_6, z30_7, z30_8, z30_9, z30_10, z30_11, z30_12, z30_13, z30_14, z30_15, z30_16, z30_17, z30_18, z30_19, z30_20, z30_21, z30_22, z30_23, z30_24, z30_25, z30_26, z30_27, z30_28, z30_29, z30_30, z30_31;
wire z31_0, z31_1, z31_2, z31_3, z31_4, z31_5, z31_6, z31_7, z31_8, z31_9, z31_10, z31_11, z31_12, z31_13, z31_14, z31_15, z31_16, z31_17, z31_18, z31_19, z31_20, z31_21, z31_22, z31_23, z31_24, z31_25, z31_26, z31_27, z31_28, z31_29, z31_30, z31_31;
wire z31_32;

wire c32 ,c33 ,c34 ,c35 ,c36 ,c37 ,c38 ,c39 ,c40 ,c41 ,c42 ,c43 ,c44 ,c45 ,c46 ,c47 ,c48 ,c49 ,c50 ,c51 ,c52 ,c53 ,c54 ,c55 ,c56 ,c57 ,c58 ,c59 ,c60 ,c61 ,c62 ,c63;
wire z32 ,z33 ,z34 ,z35 ,z36 ,z37 ,z38 ,z39 ,z40 ,z41 ,z42 ,z43 ,z44 ,z45 ,z46 ,z47 ,z48 ,z49 ,z50 ,z51 ,z52 ,z53 ,z54 ,z55 ,z56 ,z57 ,z58 ,z59 ,z60 ,z61 ,z62 ,z63;

assign X0Y0 = (X[0]&Y[0]);
assign X0Y1 = (X[0]&Y[1]);
assign X0Y2 = (X[0]&Y[2]);
assign X0Y3 = (X[0]&Y[3]);
assign X0Y4 = (X[0]&Y[4]);
assign X0Y5 = (X[0]&Y[5]);
assign X0Y6 = (X[0]&Y[6]);
assign X0Y7 = (X[0]&Y[7]);
assign X0Y8 = (X[0]&Y[8]);
assign X0Y9 = (X[0]&Y[9]);
assign X0Y10 = (X[0]&Y[10]);
assign X0Y11 = (X[0]&Y[11]);
assign X0Y12 = (X[0]&Y[12]);
assign X0Y13 = (X[0]&Y[13]);
assign X0Y14 = (X[0]&Y[14]);
assign X0Y15 = (X[0]&Y[15]);
assign X0Y16 = (X[0]&Y[16]);
assign X0Y17 = (X[0]&Y[17]);
assign X0Y18 = (X[0]&Y[18]);
assign X0Y19 = (X[0]&Y[19]);
assign X0Y20 = (X[0]&Y[20]);
assign X0Y21 = (X[0]&Y[21]);
assign X0Y22 = (X[0]&Y[22]);
assign X0Y23 = (X[0]&Y[23]);
assign X0Y24 = (X[0]&Y[24]);
assign X0Y25 = (X[0]&Y[25]);
assign X0Y26 = (X[0]&Y[26]);
assign X0Y27 = (X[0]&Y[27]);
assign X0Y28 = (X[0]&Y[28]);
assign X0Y29 = (X[0]&Y[29]);
assign X0Y30 = (X[0]&Y[30]);
assign X0Y31 = ~(X[0]&Y[31]);
assign X1Y0 = (X[1]&Y[0]);
assign X1Y1 = (X[1]&Y[1]);
assign X1Y2 = (X[1]&Y[2]);
assign X1Y3 = (X[1]&Y[3]);
assign X1Y4 = (X[1]&Y[4]);
assign X1Y5 = (X[1]&Y[5]);
assign X1Y6 = (X[1]&Y[6]);
assign X1Y7 = (X[1]&Y[7]);
assign X1Y8 = (X[1]&Y[8]);
assign X1Y9 = (X[1]&Y[9]);
assign X1Y10 = (X[1]&Y[10]);
assign X1Y11 = (X[1]&Y[11]);
assign X1Y12 = (X[1]&Y[12]);
assign X1Y13 = (X[1]&Y[13]);
assign X1Y14 = (X[1]&Y[14]);
assign X1Y15 = (X[1]&Y[15]);
assign X1Y16 = (X[1]&Y[16]);
assign X1Y17 = (X[1]&Y[17]);
assign X1Y18 = (X[1]&Y[18]);
assign X1Y19 = (X[1]&Y[19]);
assign X1Y20 = (X[1]&Y[20]);
assign X1Y21 = (X[1]&Y[21]);
assign X1Y22 = (X[1]&Y[22]);
assign X1Y23 = (X[1]&Y[23]);
assign X1Y24 = (X[1]&Y[24]);
assign X1Y25 = (X[1]&Y[25]);
assign X1Y26 = (X[1]&Y[26]);
assign X1Y27 = (X[1]&Y[27]);
assign X1Y28 = (X[1]&Y[28]);
assign X1Y29 = (X[1]&Y[29]);
assign X1Y30 = (X[1]&Y[30]);
assign X1Y31 = ~(X[1]&Y[31]);
assign X2Y0 = (X[2]&Y[0]);
assign X2Y1 = (X[2]&Y[1]);
assign X2Y2 = (X[2]&Y[2]);
assign X2Y3 = (X[2]&Y[3]);
assign X2Y4 = (X[2]&Y[4]);
assign X2Y5 = (X[2]&Y[5]);
assign X2Y6 = (X[2]&Y[6]);
assign X2Y7 = (X[2]&Y[7]);
assign X2Y8 = (X[2]&Y[8]);
assign X2Y9 = (X[2]&Y[9]);
assign X2Y10 = (X[2]&Y[10]);
assign X2Y11 = (X[2]&Y[11]);
assign X2Y12 = (X[2]&Y[12]);
assign X2Y13 = (X[2]&Y[13]);
assign X2Y14 = (X[2]&Y[14]);
assign X2Y15 = (X[2]&Y[15]);
assign X2Y16 = (X[2]&Y[16]);
assign X2Y17 = (X[2]&Y[17]);
assign X2Y18 = (X[2]&Y[18]);
assign X2Y19 = (X[2]&Y[19]);
assign X2Y20 = (X[2]&Y[20]);
assign X2Y21 = (X[2]&Y[21]);
assign X2Y22 = (X[2]&Y[22]);
assign X2Y23 = (X[2]&Y[23]);
assign X2Y24 = (X[2]&Y[24]);
assign X2Y25 = (X[2]&Y[25]);
assign X2Y26 = (X[2]&Y[26]);
assign X2Y27 = (X[2]&Y[27]);
assign X2Y28 = (X[2]&Y[28]);
assign X2Y29 = (X[2]&Y[29]);
assign X2Y30 = (X[2]&Y[30]);
assign X2Y31 = ~(X[2]&Y[31]);
assign X3Y0 = (X[3]&Y[0]);
assign X3Y1 = (X[3]&Y[1]);
assign X3Y2 = (X[3]&Y[2]);
assign X3Y3 = (X[3]&Y[3]);
assign X3Y4 = (X[3]&Y[4]);
assign X3Y5 = (X[3]&Y[5]);
assign X3Y6 = (X[3]&Y[6]);
assign X3Y7 = (X[3]&Y[7]);
assign X3Y8 = (X[3]&Y[8]);
assign X3Y9 = (X[3]&Y[9]);
assign X3Y10 = (X[3]&Y[10]);
assign X3Y11 = (X[3]&Y[11]);
assign X3Y12 = (X[3]&Y[12]);
assign X3Y13 = (X[3]&Y[13]);
assign X3Y14 = (X[3]&Y[14]);
assign X3Y15 = (X[3]&Y[15]);
assign X3Y16 = (X[3]&Y[16]);
assign X3Y17 = (X[3]&Y[17]);
assign X3Y18 = (X[3]&Y[18]);
assign X3Y19 = (X[3]&Y[19]);
assign X3Y20 = (X[3]&Y[20]);
assign X3Y21 = (X[3]&Y[21]);
assign X3Y22 = (X[3]&Y[22]);
assign X3Y23 = (X[3]&Y[23]);
assign X3Y24 = (X[3]&Y[24]);
assign X3Y25 = (X[3]&Y[25]);
assign X3Y26 = (X[3]&Y[26]);
assign X3Y27 = (X[3]&Y[27]);
assign X3Y28 = (X[3]&Y[28]);
assign X3Y29 = (X[3]&Y[29]);
assign X3Y30 = (X[3]&Y[30]);
assign X3Y31 = ~(X[3]&Y[31]);
assign X4Y0 = (X[4]&Y[0]);
assign X4Y1 = (X[4]&Y[1]);
assign X4Y2 = (X[4]&Y[2]);
assign X4Y3 = (X[4]&Y[3]);
assign X4Y4 = (X[4]&Y[4]);
assign X4Y5 = (X[4]&Y[5]);
assign X4Y6 = (X[4]&Y[6]);
assign X4Y7 = (X[4]&Y[7]);
assign X4Y8 = (X[4]&Y[8]);
assign X4Y9 = (X[4]&Y[9]);
assign X4Y10 = (X[4]&Y[10]);
assign X4Y11 = (X[4]&Y[11]);
assign X4Y12 = (X[4]&Y[12]);
assign X4Y13 = (X[4]&Y[13]);
assign X4Y14 = (X[4]&Y[14]);
assign X4Y15 = (X[4]&Y[15]);
assign X4Y16 = (X[4]&Y[16]);
assign X4Y17 = (X[4]&Y[17]);
assign X4Y18 = (X[4]&Y[18]);
assign X4Y19 = (X[4]&Y[19]);
assign X4Y20 = (X[4]&Y[20]);
assign X4Y21 = (X[4]&Y[21]);
assign X4Y22 = (X[4]&Y[22]);
assign X4Y23 = (X[4]&Y[23]);
assign X4Y24 = (X[4]&Y[24]);
assign X4Y25 = (X[4]&Y[25]);
assign X4Y26 = (X[4]&Y[26]);
assign X4Y27 = (X[4]&Y[27]);
assign X4Y28 = (X[4]&Y[28]);
assign X4Y29 = (X[4]&Y[29]);
assign X4Y30 = (X[4]&Y[30]);
assign X4Y31 = ~(X[4]&Y[31]);
assign X5Y0 = (X[5]&Y[0]);
assign X5Y1 = (X[5]&Y[1]);
assign X5Y2 = (X[5]&Y[2]);
assign X5Y3 = (X[5]&Y[3]);
assign X5Y4 = (X[5]&Y[4]);
assign X5Y5 = (X[5]&Y[5]);
assign X5Y6 = (X[5]&Y[6]);
assign X5Y7 = (X[5]&Y[7]);
assign X5Y8 = (X[5]&Y[8]);
assign X5Y9 = (X[5]&Y[9]);
assign X5Y10 = (X[5]&Y[10]);
assign X5Y11 = (X[5]&Y[11]);
assign X5Y12 = (X[5]&Y[12]);
assign X5Y13 = (X[5]&Y[13]);
assign X5Y14 = (X[5]&Y[14]);
assign X5Y15 = (X[5]&Y[15]);
assign X5Y16 = (X[5]&Y[16]);
assign X5Y17 = (X[5]&Y[17]);
assign X5Y18 = (X[5]&Y[18]);
assign X5Y19 = (X[5]&Y[19]);
assign X5Y20 = (X[5]&Y[20]);
assign X5Y21 = (X[5]&Y[21]);
assign X5Y22 = (X[5]&Y[22]);
assign X5Y23 = (X[5]&Y[23]);
assign X5Y24 = (X[5]&Y[24]);
assign X5Y25 = (X[5]&Y[25]);
assign X5Y26 = (X[5]&Y[26]);
assign X5Y27 = (X[5]&Y[27]);
assign X5Y28 = (X[5]&Y[28]);
assign X5Y29 = (X[5]&Y[29]);
assign X5Y30 = (X[5]&Y[30]);
assign X5Y31 = ~(X[5]&Y[31]);
assign X6Y0 = (X[6]&Y[0]);
assign X6Y1 = (X[6]&Y[1]);
assign X6Y2 = (X[6]&Y[2]);
assign X6Y3 = (X[6]&Y[3]);
assign X6Y4 = (X[6]&Y[4]);
assign X6Y5 = (X[6]&Y[5]);
assign X6Y6 = (X[6]&Y[6]);
assign X6Y7 = (X[6]&Y[7]);
assign X6Y8 = (X[6]&Y[8]);
assign X6Y9 = (X[6]&Y[9]);
assign X6Y10 = (X[6]&Y[10]);
assign X6Y11 = (X[6]&Y[11]);
assign X6Y12 = (X[6]&Y[12]);
assign X6Y13 = (X[6]&Y[13]);
assign X6Y14 = (X[6]&Y[14]);
assign X6Y15 = (X[6]&Y[15]);
assign X6Y16 = (X[6]&Y[16]);
assign X6Y17 = (X[6]&Y[17]);
assign X6Y18 = (X[6]&Y[18]);
assign X6Y19 = (X[6]&Y[19]);
assign X6Y20 = (X[6]&Y[20]);
assign X6Y21 = (X[6]&Y[21]);
assign X6Y22 = (X[6]&Y[22]);
assign X6Y23 = (X[6]&Y[23]);
assign X6Y24 = (X[6]&Y[24]);
assign X6Y25 = (X[6]&Y[25]);
assign X6Y26 = (X[6]&Y[26]);
assign X6Y27 = (X[6]&Y[27]);
assign X6Y28 = (X[6]&Y[28]);
assign X6Y29 = (X[6]&Y[29]);
assign X6Y30 = (X[6]&Y[30]);
assign X6Y31 = ~(X[6]&Y[31]);
assign X7Y0 = (X[7]&Y[0]);
assign X7Y1 = (X[7]&Y[1]);
assign X7Y2 = (X[7]&Y[2]);
assign X7Y3 = (X[7]&Y[3]);
assign X7Y4 = (X[7]&Y[4]);
assign X7Y5 = (X[7]&Y[5]);
assign X7Y6 = (X[7]&Y[6]);
assign X7Y7 = (X[7]&Y[7]);
assign X7Y8 = (X[7]&Y[8]);
assign X7Y9 = (X[7]&Y[9]);
assign X7Y10 = (X[7]&Y[10]);
assign X7Y11 = (X[7]&Y[11]);
assign X7Y12 = (X[7]&Y[12]);
assign X7Y13 = (X[7]&Y[13]);
assign X7Y14 = (X[7]&Y[14]);
assign X7Y15 = (X[7]&Y[15]);
assign X7Y16 = (X[7]&Y[16]);
assign X7Y17 = (X[7]&Y[17]);
assign X7Y18 = (X[7]&Y[18]);
assign X7Y19 = (X[7]&Y[19]);
assign X7Y20 = (X[7]&Y[20]);
assign X7Y21 = (X[7]&Y[21]);
assign X7Y22 = (X[7]&Y[22]);
assign X7Y23 = (X[7]&Y[23]);
assign X7Y24 = (X[7]&Y[24]);
assign X7Y25 = (X[7]&Y[25]);
assign X7Y26 = (X[7]&Y[26]);
assign X7Y27 = (X[7]&Y[27]);
assign X7Y28 = (X[7]&Y[28]);
assign X7Y29 = (X[7]&Y[29]);
assign X7Y30 = (X[7]&Y[30]);
assign X7Y31 = ~(X[7]&Y[31]);
assign X8Y0 = (X[8]&Y[0]);
assign X8Y1 = (X[8]&Y[1]);
assign X8Y2 = (X[8]&Y[2]);
assign X8Y3 = (X[8]&Y[3]);
assign X8Y4 = (X[8]&Y[4]);
assign X8Y5 = (X[8]&Y[5]);
assign X8Y6 = (X[8]&Y[6]);
assign X8Y7 = (X[8]&Y[7]);
assign X8Y8 = (X[8]&Y[8]);
assign X8Y9 = (X[8]&Y[9]);
assign X8Y10 = (X[8]&Y[10]);
assign X8Y11 = (X[8]&Y[11]);
assign X8Y12 = (X[8]&Y[12]);
assign X8Y13 = (X[8]&Y[13]);
assign X8Y14 = (X[8]&Y[14]);
assign X8Y15 = (X[8]&Y[15]);
assign X8Y16 = (X[8]&Y[16]);
assign X8Y17 = (X[8]&Y[17]);
assign X8Y18 = (X[8]&Y[18]);
assign X8Y19 = (X[8]&Y[19]);
assign X8Y20 = (X[8]&Y[20]);
assign X8Y21 = (X[8]&Y[21]);
assign X8Y22 = (X[8]&Y[22]);
assign X8Y23 = (X[8]&Y[23]);
assign X8Y24 = (X[8]&Y[24]);
assign X8Y25 = (X[8]&Y[25]);
assign X8Y26 = (X[8]&Y[26]);
assign X8Y27 = (X[8]&Y[27]);
assign X8Y28 = (X[8]&Y[28]);
assign X8Y29 = (X[8]&Y[29]);
assign X8Y30 = (X[8]&Y[30]);
assign X8Y31 = ~(X[8]&Y[31]);
assign X9Y0 = (X[9]&Y[0]);
assign X9Y1 = (X[9]&Y[1]);
assign X9Y2 = (X[9]&Y[2]);
assign X9Y3 = (X[9]&Y[3]);
assign X9Y4 = (X[9]&Y[4]);
assign X9Y5 = (X[9]&Y[5]);
assign X9Y6 = (X[9]&Y[6]);
assign X9Y7 = (X[9]&Y[7]);
assign X9Y8 = (X[9]&Y[8]);
assign X9Y9 = (X[9]&Y[9]);
assign X9Y10 = (X[9]&Y[10]);
assign X9Y11 = (X[9]&Y[11]);
assign X9Y12 = (X[9]&Y[12]);
assign X9Y13 = (X[9]&Y[13]);
assign X9Y14 = (X[9]&Y[14]);
assign X9Y15 = (X[9]&Y[15]);
assign X9Y16 = (X[9]&Y[16]);
assign X9Y17 = (X[9]&Y[17]);
assign X9Y18 = (X[9]&Y[18]);
assign X9Y19 = (X[9]&Y[19]);
assign X9Y20 = (X[9]&Y[20]);
assign X9Y21 = (X[9]&Y[21]);
assign X9Y22 = (X[9]&Y[22]);
assign X9Y23 = (X[9]&Y[23]);
assign X9Y24 = (X[9]&Y[24]);
assign X9Y25 = (X[9]&Y[25]);
assign X9Y26 = (X[9]&Y[26]);
assign X9Y27 = (X[9]&Y[27]);
assign X9Y28 = (X[9]&Y[28]);
assign X9Y29 = (X[9]&Y[29]);
assign X9Y30 = (X[9]&Y[30]);
assign X9Y31 = ~(X[9]&Y[31]);
assign X10Y0 = (X[10]&Y[0]);
assign X10Y1 = (X[10]&Y[1]);
assign X10Y2 = (X[10]&Y[2]);
assign X10Y3 = (X[10]&Y[3]);
assign X10Y4 = (X[10]&Y[4]);
assign X10Y5 = (X[10]&Y[5]);
assign X10Y6 = (X[10]&Y[6]);
assign X10Y7 = (X[10]&Y[7]);
assign X10Y8 = (X[10]&Y[8]);
assign X10Y9 = (X[10]&Y[9]);
assign X10Y10 = (X[10]&Y[10]);
assign X10Y11 = (X[10]&Y[11]);
assign X10Y12 = (X[10]&Y[12]);
assign X10Y13 = (X[10]&Y[13]);
assign X10Y14 = (X[10]&Y[14]);
assign X10Y15 = (X[10]&Y[15]);
assign X10Y16 = (X[10]&Y[16]);
assign X10Y17 = (X[10]&Y[17]);
assign X10Y18 = (X[10]&Y[18]);
assign X10Y19 = (X[10]&Y[19]);
assign X10Y20 = (X[10]&Y[20]);
assign X10Y21 = (X[10]&Y[21]);
assign X10Y22 = (X[10]&Y[22]);
assign X10Y23 = (X[10]&Y[23]);
assign X10Y24 = (X[10]&Y[24]);
assign X10Y25 = (X[10]&Y[25]);
assign X10Y26 = (X[10]&Y[26]);
assign X10Y27 = (X[10]&Y[27]);
assign X10Y28 = (X[10]&Y[28]);
assign X10Y29 = (X[10]&Y[29]);
assign X10Y30 = (X[10]&Y[30]);
assign X10Y31 = ~(X[10]&Y[31]);
assign X11Y0 = (X[11]&Y[0]);
assign X11Y1 = (X[11]&Y[1]);
assign X11Y2 = (X[11]&Y[2]);
assign X11Y3 = (X[11]&Y[3]);
assign X11Y4 = (X[11]&Y[4]);
assign X11Y5 = (X[11]&Y[5]);
assign X11Y6 = (X[11]&Y[6]);
assign X11Y7 = (X[11]&Y[7]);
assign X11Y8 = (X[11]&Y[8]);
assign X11Y9 = (X[11]&Y[9]);
assign X11Y10 = (X[11]&Y[10]);
assign X11Y11 = (X[11]&Y[11]);
assign X11Y12 = (X[11]&Y[12]);
assign X11Y13 = (X[11]&Y[13]);
assign X11Y14 = (X[11]&Y[14]);
assign X11Y15 = (X[11]&Y[15]);
assign X11Y16 = (X[11]&Y[16]);
assign X11Y17 = (X[11]&Y[17]);
assign X11Y18 = (X[11]&Y[18]);
assign X11Y19 = (X[11]&Y[19]);
assign X11Y20 = (X[11]&Y[20]);
assign X11Y21 = (X[11]&Y[21]);
assign X11Y22 = (X[11]&Y[22]);
assign X11Y23 = (X[11]&Y[23]);
assign X11Y24 = (X[11]&Y[24]);
assign X11Y25 = (X[11]&Y[25]);
assign X11Y26 = (X[11]&Y[26]);
assign X11Y27 = (X[11]&Y[27]);
assign X11Y28 = (X[11]&Y[28]);
assign X11Y29 = (X[11]&Y[29]);
assign X11Y30 = (X[11]&Y[30]);
assign X11Y31 = ~(X[11]&Y[31]);
assign X12Y0 = (X[12]&Y[0]);
assign X12Y1 = (X[12]&Y[1]);
assign X12Y2 = (X[12]&Y[2]);
assign X12Y3 = (X[12]&Y[3]);
assign X12Y4 = (X[12]&Y[4]);
assign X12Y5 = (X[12]&Y[5]);
assign X12Y6 = (X[12]&Y[6]);
assign X12Y7 = (X[12]&Y[7]);
assign X12Y8 = (X[12]&Y[8]);
assign X12Y9 = (X[12]&Y[9]);
assign X12Y10 = (X[12]&Y[10]);
assign X12Y11 = (X[12]&Y[11]);
assign X12Y12 = (X[12]&Y[12]);
assign X12Y13 = (X[12]&Y[13]);
assign X12Y14 = (X[12]&Y[14]);
assign X12Y15 = (X[12]&Y[15]);
assign X12Y16 = (X[12]&Y[16]);
assign X12Y17 = (X[12]&Y[17]);
assign X12Y18 = (X[12]&Y[18]);
assign X12Y19 = (X[12]&Y[19]);
assign X12Y20 = (X[12]&Y[20]);
assign X12Y21 = (X[12]&Y[21]);
assign X12Y22 = (X[12]&Y[22]);
assign X12Y23 = (X[12]&Y[23]);
assign X12Y24 = (X[12]&Y[24]);
assign X12Y25 = (X[12]&Y[25]);
assign X12Y26 = (X[12]&Y[26]);
assign X12Y27 = (X[12]&Y[27]);
assign X12Y28 = (X[12]&Y[28]);
assign X12Y29 = (X[12]&Y[29]);
assign X12Y30 = (X[12]&Y[30]);
assign X12Y31 = ~(X[12]&Y[31]);
assign X13Y0 = (X[13]&Y[0]);
assign X13Y1 = (X[13]&Y[1]);
assign X13Y2 = (X[13]&Y[2]);
assign X13Y3 = (X[13]&Y[3]);
assign X13Y4 = (X[13]&Y[4]);
assign X13Y5 = (X[13]&Y[5]);
assign X13Y6 = (X[13]&Y[6]);
assign X13Y7 = (X[13]&Y[7]);
assign X13Y8 = (X[13]&Y[8]);
assign X13Y9 = (X[13]&Y[9]);
assign X13Y10 = (X[13]&Y[10]);
assign X13Y11 = (X[13]&Y[11]);
assign X13Y12 = (X[13]&Y[12]);
assign X13Y13 = (X[13]&Y[13]);
assign X13Y14 = (X[13]&Y[14]);
assign X13Y15 = (X[13]&Y[15]);
assign X13Y16 = (X[13]&Y[16]);
assign X13Y17 = (X[13]&Y[17]);
assign X13Y18 = (X[13]&Y[18]);
assign X13Y19 = (X[13]&Y[19]);
assign X13Y20 = (X[13]&Y[20]);
assign X13Y21 = (X[13]&Y[21]);
assign X13Y22 = (X[13]&Y[22]);
assign X13Y23 = (X[13]&Y[23]);
assign X13Y24 = (X[13]&Y[24]);
assign X13Y25 = (X[13]&Y[25]);
assign X13Y26 = (X[13]&Y[26]);
assign X13Y27 = (X[13]&Y[27]);
assign X13Y28 = (X[13]&Y[28]);
assign X13Y29 = (X[13]&Y[29]);
assign X13Y30 = (X[13]&Y[30]);
assign X13Y31 = ~(X[13]&Y[31]);
assign X14Y0 = (X[14]&Y[0]);
assign X14Y1 = (X[14]&Y[1]);
assign X14Y2 = (X[14]&Y[2]);
assign X14Y3 = (X[14]&Y[3]);
assign X14Y4 = (X[14]&Y[4]);
assign X14Y5 = (X[14]&Y[5]);
assign X14Y6 = (X[14]&Y[6]);
assign X14Y7 = (X[14]&Y[7]);
assign X14Y8 = (X[14]&Y[8]);
assign X14Y9 = (X[14]&Y[9]);
assign X14Y10 = (X[14]&Y[10]);
assign X14Y11 = (X[14]&Y[11]);
assign X14Y12 = (X[14]&Y[12]);
assign X14Y13 = (X[14]&Y[13]);
assign X14Y14 = (X[14]&Y[14]);
assign X14Y15 = (X[14]&Y[15]);
assign X14Y16 = (X[14]&Y[16]);
assign X14Y17 = (X[14]&Y[17]);
assign X14Y18 = (X[14]&Y[18]);
assign X14Y19 = (X[14]&Y[19]);
assign X14Y20 = (X[14]&Y[20]);
assign X14Y21 = (X[14]&Y[21]);
assign X14Y22 = (X[14]&Y[22]);
assign X14Y23 = (X[14]&Y[23]);
assign X14Y24 = (X[14]&Y[24]);
assign X14Y25 = (X[14]&Y[25]);
assign X14Y26 = (X[14]&Y[26]);
assign X14Y27 = (X[14]&Y[27]);
assign X14Y28 = (X[14]&Y[28]);
assign X14Y29 = (X[14]&Y[29]);
assign X14Y30 = (X[14]&Y[30]);
assign X14Y31 = ~(X[14]&Y[31]);
assign X15Y0 = (X[15]&Y[0]);
assign X15Y1 = (X[15]&Y[1]);
assign X15Y2 = (X[15]&Y[2]);
assign X15Y3 = (X[15]&Y[3]);
assign X15Y4 = (X[15]&Y[4]);
assign X15Y5 = (X[15]&Y[5]);
assign X15Y6 = (X[15]&Y[6]);
assign X15Y7 = (X[15]&Y[7]);
assign X15Y8 = (X[15]&Y[8]);
assign X15Y9 = (X[15]&Y[9]);
assign X15Y10 = (X[15]&Y[10]);
assign X15Y11 = (X[15]&Y[11]);
assign X15Y12 = (X[15]&Y[12]);
assign X15Y13 = (X[15]&Y[13]);
assign X15Y14 = (X[15]&Y[14]);
assign X15Y15 = (X[15]&Y[15]);
assign X15Y16 = (X[15]&Y[16]);
assign X15Y17 = (X[15]&Y[17]);
assign X15Y18 = (X[15]&Y[18]);
assign X15Y19 = (X[15]&Y[19]);
assign X15Y20 = (X[15]&Y[20]);
assign X15Y21 = (X[15]&Y[21]);
assign X15Y22 = (X[15]&Y[22]);
assign X15Y23 = (X[15]&Y[23]);
assign X15Y24 = (X[15]&Y[24]);
assign X15Y25 = (X[15]&Y[25]);
assign X15Y26 = (X[15]&Y[26]);
assign X15Y27 = (X[15]&Y[27]);
assign X15Y28 = (X[15]&Y[28]);
assign X15Y29 = (X[15]&Y[29]);
assign X15Y30 = (X[15]&Y[30]);
assign X15Y31 = ~(X[15]&Y[31]);
assign X16Y0 = (X[16]&Y[0]);
assign X16Y1 = (X[16]&Y[1]);
assign X16Y2 = (X[16]&Y[2]);
assign X16Y3 = (X[16]&Y[3]);
assign X16Y4 = (X[16]&Y[4]);
assign X16Y5 = (X[16]&Y[5]);
assign X16Y6 = (X[16]&Y[6]);
assign X16Y7 = (X[16]&Y[7]);
assign X16Y8 = (X[16]&Y[8]);
assign X16Y9 = (X[16]&Y[9]);
assign X16Y10 = (X[16]&Y[10]);
assign X16Y11 = (X[16]&Y[11]);
assign X16Y12 = (X[16]&Y[12]);
assign X16Y13 = (X[16]&Y[13]);
assign X16Y14 = (X[16]&Y[14]);
assign X16Y15 = (X[16]&Y[15]);
assign X16Y16 = (X[16]&Y[16]);
assign X16Y17 = (X[16]&Y[17]);
assign X16Y18 = (X[16]&Y[18]);
assign X16Y19 = (X[16]&Y[19]);
assign X16Y20 = (X[16]&Y[20]);
assign X16Y21 = (X[16]&Y[21]);
assign X16Y22 = (X[16]&Y[22]);
assign X16Y23 = (X[16]&Y[23]);
assign X16Y24 = (X[16]&Y[24]);
assign X16Y25 = (X[16]&Y[25]);
assign X16Y26 = (X[16]&Y[26]);
assign X16Y27 = (X[16]&Y[27]);
assign X16Y28 = (X[16]&Y[28]);
assign X16Y29 = (X[16]&Y[29]);
assign X16Y30 = (X[16]&Y[30]);
assign X16Y31 = ~(X[16]&Y[31]);
assign X17Y0 = (X[17]&Y[0]);
assign X17Y1 = (X[17]&Y[1]);
assign X17Y2 = (X[17]&Y[2]);
assign X17Y3 = (X[17]&Y[3]);
assign X17Y4 = (X[17]&Y[4]);
assign X17Y5 = (X[17]&Y[5]);
assign X17Y6 = (X[17]&Y[6]);
assign X17Y7 = (X[17]&Y[7]);
assign X17Y8 = (X[17]&Y[8]);
assign X17Y9 = (X[17]&Y[9]);
assign X17Y10 = (X[17]&Y[10]);
assign X17Y11 = (X[17]&Y[11]);
assign X17Y12 = (X[17]&Y[12]);
assign X17Y13 = (X[17]&Y[13]);
assign X17Y14 = (X[17]&Y[14]);
assign X17Y15 = (X[17]&Y[15]);
assign X17Y16 = (X[17]&Y[16]);
assign X17Y17 = (X[17]&Y[17]);
assign X17Y18 = (X[17]&Y[18]);
assign X17Y19 = (X[17]&Y[19]);
assign X17Y20 = (X[17]&Y[20]);
assign X17Y21 = (X[17]&Y[21]);
assign X17Y22 = (X[17]&Y[22]);
assign X17Y23 = (X[17]&Y[23]);
assign X17Y24 = (X[17]&Y[24]);
assign X17Y25 = (X[17]&Y[25]);
assign X17Y26 = (X[17]&Y[26]);
assign X17Y27 = (X[17]&Y[27]);
assign X17Y28 = (X[17]&Y[28]);
assign X17Y29 = (X[17]&Y[29]);
assign X17Y30 = (X[17]&Y[30]);
assign X17Y31 = ~(X[17]&Y[31]);
assign X18Y0 = (X[18]&Y[0]);
assign X18Y1 = (X[18]&Y[1]);
assign X18Y2 = (X[18]&Y[2]);
assign X18Y3 = (X[18]&Y[3]);
assign X18Y4 = (X[18]&Y[4]);
assign X18Y5 = (X[18]&Y[5]);
assign X18Y6 = (X[18]&Y[6]);
assign X18Y7 = (X[18]&Y[7]);
assign X18Y8 = (X[18]&Y[8]);
assign X18Y9 = (X[18]&Y[9]);
assign X18Y10 = (X[18]&Y[10]);
assign X18Y11 = (X[18]&Y[11]);
assign X18Y12 = (X[18]&Y[12]);
assign X18Y13 = (X[18]&Y[13]);
assign X18Y14 = (X[18]&Y[14]);
assign X18Y15 = (X[18]&Y[15]);
assign X18Y16 = (X[18]&Y[16]);
assign X18Y17 = (X[18]&Y[17]);
assign X18Y18 = (X[18]&Y[18]);
assign X18Y19 = (X[18]&Y[19]);
assign X18Y20 = (X[18]&Y[20]);
assign X18Y21 = (X[18]&Y[21]);
assign X18Y22 = (X[18]&Y[22]);
assign X18Y23 = (X[18]&Y[23]);
assign X18Y24 = (X[18]&Y[24]);
assign X18Y25 = (X[18]&Y[25]);
assign X18Y26 = (X[18]&Y[26]);
assign X18Y27 = (X[18]&Y[27]);
assign X18Y28 = (X[18]&Y[28]);
assign X18Y29 = (X[18]&Y[29]);
assign X18Y30 = (X[18]&Y[30]);
assign X18Y31 = ~(X[18]&Y[31]);
assign X19Y0 = (X[19]&Y[0]);
assign X19Y1 = (X[19]&Y[1]);
assign X19Y2 = (X[19]&Y[2]);
assign X19Y3 = (X[19]&Y[3]);
assign X19Y4 = (X[19]&Y[4]);
assign X19Y5 = (X[19]&Y[5]);
assign X19Y6 = (X[19]&Y[6]);
assign X19Y7 = (X[19]&Y[7]);
assign X19Y8 = (X[19]&Y[8]);
assign X19Y9 = (X[19]&Y[9]);
assign X19Y10 = (X[19]&Y[10]);
assign X19Y11 = (X[19]&Y[11]);
assign X19Y12 = (X[19]&Y[12]);
assign X19Y13 = (X[19]&Y[13]);
assign X19Y14 = (X[19]&Y[14]);
assign X19Y15 = (X[19]&Y[15]);
assign X19Y16 = (X[19]&Y[16]);
assign X19Y17 = (X[19]&Y[17]);
assign X19Y18 = (X[19]&Y[18]);
assign X19Y19 = (X[19]&Y[19]);
assign X19Y20 = (X[19]&Y[20]);
assign X19Y21 = (X[19]&Y[21]);
assign X19Y22 = (X[19]&Y[22]);
assign X19Y23 = (X[19]&Y[23]);
assign X19Y24 = (X[19]&Y[24]);
assign X19Y25 = (X[19]&Y[25]);
assign X19Y26 = (X[19]&Y[26]);
assign X19Y27 = (X[19]&Y[27]);
assign X19Y28 = (X[19]&Y[28]);
assign X19Y29 = (X[19]&Y[29]);
assign X19Y30 = (X[19]&Y[30]);
assign X19Y31 = ~(X[19]&Y[31]);
assign X20Y0 = (X[20]&Y[0]);
assign X20Y1 = (X[20]&Y[1]);
assign X20Y2 = (X[20]&Y[2]);
assign X20Y3 = (X[20]&Y[3]);
assign X20Y4 = (X[20]&Y[4]);
assign X20Y5 = (X[20]&Y[5]);
assign X20Y6 = (X[20]&Y[6]);
assign X20Y7 = (X[20]&Y[7]);
assign X20Y8 = (X[20]&Y[8]);
assign X20Y9 = (X[20]&Y[9]);
assign X20Y10 = (X[20]&Y[10]);
assign X20Y11 = (X[20]&Y[11]);
assign X20Y12 = (X[20]&Y[12]);
assign X20Y13 = (X[20]&Y[13]);
assign X20Y14 = (X[20]&Y[14]);
assign X20Y15 = (X[20]&Y[15]);
assign X20Y16 = (X[20]&Y[16]);
assign X20Y17 = (X[20]&Y[17]);
assign X20Y18 = (X[20]&Y[18]);
assign X20Y19 = (X[20]&Y[19]);
assign X20Y20 = (X[20]&Y[20]);
assign X20Y21 = (X[20]&Y[21]);
assign X20Y22 = (X[20]&Y[22]);
assign X20Y23 = (X[20]&Y[23]);
assign X20Y24 = (X[20]&Y[24]);
assign X20Y25 = (X[20]&Y[25]);
assign X20Y26 = (X[20]&Y[26]);
assign X20Y27 = (X[20]&Y[27]);
assign X20Y28 = (X[20]&Y[28]);
assign X20Y29 = (X[20]&Y[29]);
assign X20Y30 = (X[20]&Y[30]);
assign X20Y31 = ~(X[20]&Y[31]);
assign X21Y0 = (X[21]&Y[0]);
assign X21Y1 = (X[21]&Y[1]);
assign X21Y2 = (X[21]&Y[2]);
assign X21Y3 = (X[21]&Y[3]);
assign X21Y4 = (X[21]&Y[4]);
assign X21Y5 = (X[21]&Y[5]);
assign X21Y6 = (X[21]&Y[6]);
assign X21Y7 = (X[21]&Y[7]);
assign X21Y8 = (X[21]&Y[8]);
assign X21Y9 = (X[21]&Y[9]);
assign X21Y10 = (X[21]&Y[10]);
assign X21Y11 = (X[21]&Y[11]);
assign X21Y12 = (X[21]&Y[12]);
assign X21Y13 = (X[21]&Y[13]);
assign X21Y14 = (X[21]&Y[14]);
assign X21Y15 = (X[21]&Y[15]);
assign X21Y16 = (X[21]&Y[16]);
assign X21Y17 = (X[21]&Y[17]);
assign X21Y18 = (X[21]&Y[18]);
assign X21Y19 = (X[21]&Y[19]);
assign X21Y20 = (X[21]&Y[20]);
assign X21Y21 = (X[21]&Y[21]);
assign X21Y22 = (X[21]&Y[22]);
assign X21Y23 = (X[21]&Y[23]);
assign X21Y24 = (X[21]&Y[24]);
assign X21Y25 = (X[21]&Y[25]);
assign X21Y26 = (X[21]&Y[26]);
assign X21Y27 = (X[21]&Y[27]);
assign X21Y28 = (X[21]&Y[28]);
assign X21Y29 = (X[21]&Y[29]);
assign X21Y30 = (X[21]&Y[30]);
assign X21Y31 = ~(X[21]&Y[31]);
assign X22Y0 = (X[22]&Y[0]);
assign X22Y1 = (X[22]&Y[1]);
assign X22Y2 = (X[22]&Y[2]);
assign X22Y3 = (X[22]&Y[3]);
assign X22Y4 = (X[22]&Y[4]);
assign X22Y5 = (X[22]&Y[5]);
assign X22Y6 = (X[22]&Y[6]);
assign X22Y7 = (X[22]&Y[7]);
assign X22Y8 = (X[22]&Y[8]);
assign X22Y9 = (X[22]&Y[9]);
assign X22Y10 = (X[22]&Y[10]);
assign X22Y11 = (X[22]&Y[11]);
assign X22Y12 = (X[22]&Y[12]);
assign X22Y13 = (X[22]&Y[13]);
assign X22Y14 = (X[22]&Y[14]);
assign X22Y15 = (X[22]&Y[15]);
assign X22Y16 = (X[22]&Y[16]);
assign X22Y17 = (X[22]&Y[17]);
assign X22Y18 = (X[22]&Y[18]);
assign X22Y19 = (X[22]&Y[19]);
assign X22Y20 = (X[22]&Y[20]);
assign X22Y21 = (X[22]&Y[21]);
assign X22Y22 = (X[22]&Y[22]);
assign X22Y23 = (X[22]&Y[23]);
assign X22Y24 = (X[22]&Y[24]);
assign X22Y25 = (X[22]&Y[25]);
assign X22Y26 = (X[22]&Y[26]);
assign X22Y27 = (X[22]&Y[27]);
assign X22Y28 = (X[22]&Y[28]);
assign X22Y29 = (X[22]&Y[29]);
assign X22Y30 = (X[22]&Y[30]);
assign X22Y31 = ~(X[22]&Y[31]);
assign X23Y0 = (X[23]&Y[0]);
assign X23Y1 = (X[23]&Y[1]);
assign X23Y2 = (X[23]&Y[2]);
assign X23Y3 = (X[23]&Y[3]);
assign X23Y4 = (X[23]&Y[4]);
assign X23Y5 = (X[23]&Y[5]);
assign X23Y6 = (X[23]&Y[6]);
assign X23Y7 = (X[23]&Y[7]);
assign X23Y8 = (X[23]&Y[8]);
assign X23Y9 = (X[23]&Y[9]);
assign X23Y10 = (X[23]&Y[10]);
assign X23Y11 = (X[23]&Y[11]);
assign X23Y12 = (X[23]&Y[12]);
assign X23Y13 = (X[23]&Y[13]);
assign X23Y14 = (X[23]&Y[14]);
assign X23Y15 = (X[23]&Y[15]);
assign X23Y16 = (X[23]&Y[16]);
assign X23Y17 = (X[23]&Y[17]);
assign X23Y18 = (X[23]&Y[18]);
assign X23Y19 = (X[23]&Y[19]);
assign X23Y20 = (X[23]&Y[20]);
assign X23Y21 = (X[23]&Y[21]);
assign X23Y22 = (X[23]&Y[22]);
assign X23Y23 = (X[23]&Y[23]);
assign X23Y24 = (X[23]&Y[24]);
assign X23Y25 = (X[23]&Y[25]);
assign X23Y26 = (X[23]&Y[26]);
assign X23Y27 = (X[23]&Y[27]);
assign X23Y28 = (X[23]&Y[28]);
assign X23Y29 = (X[23]&Y[29]);
assign X23Y30 = (X[23]&Y[30]);
assign X23Y31 = ~(X[23]&Y[31]);
assign X24Y0 = (X[24]&Y[0]);
assign X24Y1 = (X[24]&Y[1]);
assign X24Y2 = (X[24]&Y[2]);
assign X24Y3 = (X[24]&Y[3]);
assign X24Y4 = (X[24]&Y[4]);
assign X24Y5 = (X[24]&Y[5]);
assign X24Y6 = (X[24]&Y[6]);
assign X24Y7 = (X[24]&Y[7]);
assign X24Y8 = (X[24]&Y[8]);
assign X24Y9 = (X[24]&Y[9]);
assign X24Y10 = (X[24]&Y[10]);
assign X24Y11 = (X[24]&Y[11]);
assign X24Y12 = (X[24]&Y[12]);
assign X24Y13 = (X[24]&Y[13]);
assign X24Y14 = (X[24]&Y[14]);
assign X24Y15 = (X[24]&Y[15]);
assign X24Y16 = (X[24]&Y[16]);
assign X24Y17 = (X[24]&Y[17]);
assign X24Y18 = (X[24]&Y[18]);
assign X24Y19 = (X[24]&Y[19]);
assign X24Y20 = (X[24]&Y[20]);
assign X24Y21 = (X[24]&Y[21]);
assign X24Y22 = (X[24]&Y[22]);
assign X24Y23 = (X[24]&Y[23]);
assign X24Y24 = (X[24]&Y[24]);
assign X24Y25 = (X[24]&Y[25]);
assign X24Y26 = (X[24]&Y[26]);
assign X24Y27 = (X[24]&Y[27]);
assign X24Y28 = (X[24]&Y[28]);
assign X24Y29 = (X[24]&Y[29]);
assign X24Y30 = (X[24]&Y[30]);
assign X24Y31 = ~(X[24]&Y[31]);
assign X25Y0 = (X[25]&Y[0]);
assign X25Y1 = (X[25]&Y[1]);
assign X25Y2 = (X[25]&Y[2]);
assign X25Y3 = (X[25]&Y[3]);
assign X25Y4 = (X[25]&Y[4]);
assign X25Y5 = (X[25]&Y[5]);
assign X25Y6 = (X[25]&Y[6]);
assign X25Y7 = (X[25]&Y[7]);
assign X25Y8 = (X[25]&Y[8]);
assign X25Y9 = (X[25]&Y[9]);
assign X25Y10 = (X[25]&Y[10]);
assign X25Y11 = (X[25]&Y[11]);
assign X25Y12 = (X[25]&Y[12]);
assign X25Y13 = (X[25]&Y[13]);
assign X25Y14 = (X[25]&Y[14]);
assign X25Y15 = (X[25]&Y[15]);
assign X25Y16 = (X[25]&Y[16]);
assign X25Y17 = (X[25]&Y[17]);
assign X25Y18 = (X[25]&Y[18]);
assign X25Y19 = (X[25]&Y[19]);
assign X25Y20 = (X[25]&Y[20]);
assign X25Y21 = (X[25]&Y[21]);
assign X25Y22 = (X[25]&Y[22]);
assign X25Y23 = (X[25]&Y[23]);
assign X25Y24 = (X[25]&Y[24]);
assign X25Y25 = (X[25]&Y[25]);
assign X25Y26 = (X[25]&Y[26]);
assign X25Y27 = (X[25]&Y[27]);
assign X25Y28 = (X[25]&Y[28]);
assign X25Y29 = (X[25]&Y[29]);
assign X25Y30 = (X[25]&Y[30]);
assign X25Y31 = ~(X[25]&Y[31]);
assign X26Y0 = (X[26]&Y[0]);
assign X26Y1 = (X[26]&Y[1]);
assign X26Y2 = (X[26]&Y[2]);
assign X26Y3 = (X[26]&Y[3]);
assign X26Y4 = (X[26]&Y[4]);
assign X26Y5 = (X[26]&Y[5]);
assign X26Y6 = (X[26]&Y[6]);
assign X26Y7 = (X[26]&Y[7]);
assign X26Y8 = (X[26]&Y[8]);
assign X26Y9 = (X[26]&Y[9]);
assign X26Y10 = (X[26]&Y[10]);
assign X26Y11 = (X[26]&Y[11]);
assign X26Y12 = (X[26]&Y[12]);
assign X26Y13 = (X[26]&Y[13]);
assign X26Y14 = (X[26]&Y[14]);
assign X26Y15 = (X[26]&Y[15]);
assign X26Y16 = (X[26]&Y[16]);
assign X26Y17 = (X[26]&Y[17]);
assign X26Y18 = (X[26]&Y[18]);
assign X26Y19 = (X[26]&Y[19]);
assign X26Y20 = (X[26]&Y[20]);
assign X26Y21 = (X[26]&Y[21]);
assign X26Y22 = (X[26]&Y[22]);
assign X26Y23 = (X[26]&Y[23]);
assign X26Y24 = (X[26]&Y[24]);
assign X26Y25 = (X[26]&Y[25]);
assign X26Y26 = (X[26]&Y[26]);
assign X26Y27 = (X[26]&Y[27]);
assign X26Y28 = (X[26]&Y[28]);
assign X26Y29 = (X[26]&Y[29]);
assign X26Y30 = (X[26]&Y[30]);
assign X26Y31 = ~(X[26]&Y[31]);
assign X27Y0 = (X[27]&Y[0]);
assign X27Y1 = (X[27]&Y[1]);
assign X27Y2 = (X[27]&Y[2]);
assign X27Y3 = (X[27]&Y[3]);
assign X27Y4 = (X[27]&Y[4]);
assign X27Y5 = (X[27]&Y[5]);
assign X27Y6 = (X[27]&Y[6]);
assign X27Y7 = (X[27]&Y[7]);
assign X27Y8 = (X[27]&Y[8]);
assign X27Y9 = (X[27]&Y[9]);
assign X27Y10 = (X[27]&Y[10]);
assign X27Y11 = (X[27]&Y[11]);
assign X27Y12 = (X[27]&Y[12]);
assign X27Y13 = (X[27]&Y[13]);
assign X27Y14 = (X[27]&Y[14]);
assign X27Y15 = (X[27]&Y[15]);
assign X27Y16 = (X[27]&Y[16]);
assign X27Y17 = (X[27]&Y[17]);
assign X27Y18 = (X[27]&Y[18]);
assign X27Y19 = (X[27]&Y[19]);
assign X27Y20 = (X[27]&Y[20]);
assign X27Y21 = (X[27]&Y[21]);
assign X27Y22 = (X[27]&Y[22]);
assign X27Y23 = (X[27]&Y[23]);
assign X27Y24 = (X[27]&Y[24]);
assign X27Y25 = (X[27]&Y[25]);
assign X27Y26 = (X[27]&Y[26]);
assign X27Y27 = (X[27]&Y[27]);
assign X27Y28 = (X[27]&Y[28]);
assign X27Y29 = (X[27]&Y[29]);
assign X27Y30 = (X[27]&Y[30]);
assign X27Y31 = ~(X[27]&Y[31]);
assign X28Y0 = (X[28]&Y[0]);
assign X28Y1 = (X[28]&Y[1]);
assign X28Y2 = (X[28]&Y[2]);
assign X28Y3 = (X[28]&Y[3]);
assign X28Y4 = (X[28]&Y[4]);
assign X28Y5 = (X[28]&Y[5]);
assign X28Y6 = (X[28]&Y[6]);
assign X28Y7 = (X[28]&Y[7]);
assign X28Y8 = (X[28]&Y[8]);
assign X28Y9 = (X[28]&Y[9]);
assign X28Y10 = (X[28]&Y[10]);
assign X28Y11 = (X[28]&Y[11]);
assign X28Y12 = (X[28]&Y[12]);
assign X28Y13 = (X[28]&Y[13]);
assign X28Y14 = (X[28]&Y[14]);
assign X28Y15 = (X[28]&Y[15]);
assign X28Y16 = (X[28]&Y[16]);
assign X28Y17 = (X[28]&Y[17]);
assign X28Y18 = (X[28]&Y[18]);
assign X28Y19 = (X[28]&Y[19]);
assign X28Y20 = (X[28]&Y[20]);
assign X28Y21 = (X[28]&Y[21]);
assign X28Y22 = (X[28]&Y[22]);
assign X28Y23 = (X[28]&Y[23]);
assign X28Y24 = (X[28]&Y[24]);
assign X28Y25 = (X[28]&Y[25]);
assign X28Y26 = (X[28]&Y[26]);
assign X28Y27 = (X[28]&Y[27]);
assign X28Y28 = (X[28]&Y[28]);
assign X28Y29 = (X[28]&Y[29]);
assign X28Y30 = (X[28]&Y[30]);
assign X28Y31 = ~(X[28]&Y[31]);
assign X29Y0 = (X[29]&Y[0]);
assign X29Y1 = (X[29]&Y[1]);
assign X29Y2 = (X[29]&Y[2]);
assign X29Y3 = (X[29]&Y[3]);
assign X29Y4 = (X[29]&Y[4]);
assign X29Y5 = (X[29]&Y[5]);
assign X29Y6 = (X[29]&Y[6]);
assign X29Y7 = (X[29]&Y[7]);
assign X29Y8 = (X[29]&Y[8]);
assign X29Y9 = (X[29]&Y[9]);
assign X29Y10 = (X[29]&Y[10]);
assign X29Y11 = (X[29]&Y[11]);
assign X29Y12 = (X[29]&Y[12]);
assign X29Y13 = (X[29]&Y[13]);
assign X29Y14 = (X[29]&Y[14]);
assign X29Y15 = (X[29]&Y[15]);
assign X29Y16 = (X[29]&Y[16]);
assign X29Y17 = (X[29]&Y[17]);
assign X29Y18 = (X[29]&Y[18]);
assign X29Y19 = (X[29]&Y[19]);
assign X29Y20 = (X[29]&Y[20]);
assign X29Y21 = (X[29]&Y[21]);
assign X29Y22 = (X[29]&Y[22]);
assign X29Y23 = (X[29]&Y[23]);
assign X29Y24 = (X[29]&Y[24]);
assign X29Y25 = (X[29]&Y[25]);
assign X29Y26 = (X[29]&Y[26]);
assign X29Y27 = (X[29]&Y[27]);
assign X29Y28 = (X[29]&Y[28]);
assign X29Y29 = (X[29]&Y[29]);
assign X29Y30 = (X[29]&Y[30]);
assign X29Y31 = ~(X[29]&Y[31]);
assign X30Y0 = (X[30]&Y[0]);
assign X30Y1 = (X[30]&Y[1]);
assign X30Y2 = (X[30]&Y[2]);
assign X30Y3 = (X[30]&Y[3]);
assign X30Y4 = (X[30]&Y[4]);
assign X30Y5 = (X[30]&Y[5]);
assign X30Y6 = (X[30]&Y[6]);
assign X30Y7 = (X[30]&Y[7]);
assign X30Y8 = (X[30]&Y[8]);
assign X30Y9 = (X[30]&Y[9]);
assign X30Y10 = (X[30]&Y[10]);
assign X30Y11 = (X[30]&Y[11]);
assign X30Y12 = (X[30]&Y[12]);
assign X30Y13 = (X[30]&Y[13]);
assign X30Y14 = (X[30]&Y[14]);
assign X30Y15 = (X[30]&Y[15]);
assign X30Y16 = (X[30]&Y[16]);
assign X30Y17 = (X[30]&Y[17]);
assign X30Y18 = (X[30]&Y[18]);
assign X30Y19 = (X[30]&Y[19]);
assign X30Y20 = (X[30]&Y[20]);
assign X30Y21 = (X[30]&Y[21]);
assign X30Y22 = (X[30]&Y[22]);
assign X30Y23 = (X[30]&Y[23]);
assign X30Y24 = (X[30]&Y[24]);
assign X30Y25 = (X[30]&Y[25]);
assign X30Y26 = (X[30]&Y[26]);
assign X30Y27 = (X[30]&Y[27]);
assign X30Y28 = (X[30]&Y[28]);
assign X30Y29 = (X[30]&Y[29]);
assign X30Y30 = (X[30]&Y[30]);
assign X30Y31 = ~(X[30]&Y[31]);
assign X31Y0 = ~(X[31]&Y[0]);
assign X31Y1 = ~(X[31]&Y[1]);
assign X31Y2 = ~(X[31]&Y[2]);
assign X31Y3 = ~(X[31]&Y[3]);
assign X31Y4 = ~(X[31]&Y[4]);
assign X31Y5 = ~(X[31]&Y[5]);
assign X31Y6 = ~(X[31]&Y[6]);
assign X31Y7 = ~(X[31]&Y[7]);
assign X31Y8 = ~(X[31]&Y[8]);
assign X31Y9 = ~(X[31]&Y[9]);
assign X31Y10 = ~(X[31]&Y[10]);
assign X31Y11 = ~(X[31]&Y[11]);
assign X31Y12 = ~(X[31]&Y[12]);
assign X31Y13 = ~(X[31]&Y[13]);
assign X31Y14 = ~(X[31]&Y[14]);
assign X31Y15 = ~(X[31]&Y[15]);
assign X31Y16 = ~(X[31]&Y[16]);
assign X31Y17 = ~(X[31]&Y[17]);
assign X31Y18 = ~(X[31]&Y[18]);
assign X31Y19 = ~(X[31]&Y[19]);
assign X31Y20 = ~(X[31]&Y[20]);
assign X31Y21 = ~(X[31]&Y[21]);
assign X31Y22 = ~(X[31]&Y[22]);
assign X31Y23 = ~(X[31]&Y[23]);
assign X31Y24 = ~(X[31]&Y[24]);
assign X31Y25 = ~(X[31]&Y[25]);
assign X31Y26 = ~(X[31]&Y[26]);
assign X31Y27 = ~(X[31]&Y[27]);
assign X31Y28 = ~(X[31]&Y[28]);
assign X31Y29 = ~(X[31]&Y[29]);
assign X31Y30 = ~(X[31]&Y[30]);
assign X31Y31 = (X[31]&Y[31]);

assign c0_31 = 1;
HA h1_0(X0Y1,X1Y0,c1_0,z1_0);
HA h1_1(X1Y1,X2Y0,c1_1,z1_1);
HA h1_2(X2Y1,X3Y0,c1_2,z1_2);
HA h1_3(X3Y1,X4Y0,c1_3,z1_3);
HA h1_4(X4Y1,X5Y0,c1_4,z1_4);
HA h1_5(X5Y1,X6Y0,c1_5,z1_5);
HA h1_6(X6Y1,X7Y0,c1_6,z1_6);
HA h1_7(X7Y1,X8Y0,c1_7,z1_7);
HA h1_8(X8Y1,X9Y0,c1_8,z1_8);
HA h1_9(X9Y1,X10Y0,c1_9,z1_9);
HA h1_10(X10Y1,X11Y0,c1_10,z1_10);
HA h1_11(X11Y1,X12Y0,c1_11,z1_11);
HA h1_12(X12Y1,X13Y0,c1_12,z1_12);
HA h1_13(X13Y1,X14Y0,c1_13,z1_13);
HA h1_14(X14Y1,X15Y0,c1_14,z1_14);
HA h1_15(X15Y1,X16Y0,c1_15,z1_15);
HA h1_16(X16Y1,X17Y0,c1_16,z1_16);
HA h1_17(X17Y1,X18Y0,c1_17,z1_17);
HA h1_18(X18Y1,X19Y0,c1_18,z1_18);
HA h1_19(X19Y1,X20Y0,c1_19,z1_19);
HA h1_20(X20Y1,X21Y0,c1_20,z1_20);
HA h1_21(X21Y1,X22Y0,c1_21,z1_21);
HA h1_22(X22Y1,X23Y0,c1_22,z1_22);
HA h1_23(X23Y1,X24Y0,c1_23,z1_23);
HA h1_24(X24Y1,X25Y0,c1_24,z1_24);
HA h1_25(X25Y1,X26Y0,c1_25,z1_25);
HA h1_26(X26Y1,X27Y0,c1_26,z1_26);
HA h1_27(X27Y1,X28Y0,c1_27,z1_27);
HA h1_28(X28Y1,X29Y0,c1_28,z1_28);
HA h1_29(X29Y1,X30Y0,c1_29,z1_29);
HA h1_30(X30Y1,X31Y0,c1_30,z1_30);
HA h1_31(X31Y1,c0_31,c1_31,z1_31);
HA h2_31(X31Y2,c1_31,c2_31,z2_31);
HA h3_31(X31Y3,c2_31,c3_31,z3_31);
HA h4_31(X31Y4,c3_31,c4_31,z4_31);
HA h5_31(X31Y5,c4_31,c5_31,z5_31);
HA h6_31(X31Y6,c5_31,c6_31,z6_31);
HA h7_31(X31Y7,c6_31,c7_31,z7_31);
HA h8_31(X31Y8,c7_31,c8_31,z8_31);
HA h9_31(X31Y9,c8_31,c9_31,z9_31);
HA h10_31(X31Y10,c9_31,c10_31,z10_31);
HA h11_31(X31Y11,c10_31,c11_31,z11_31);
HA h12_31(X31Y12,c11_31,c12_31,z12_31);
HA h13_31(X31Y13,c12_31,c13_31,z13_31);
HA h14_31(X31Y14,c13_31,c14_31,z14_31);
HA h15_31(X31Y15,c14_31,c15_31,z15_31);
HA h16_31(X31Y16,c15_31,c16_31,z16_31);
HA h17_31(X31Y17,c16_31,c17_31,z17_31);
HA h18_31(X31Y18,c17_31,c18_31,z18_31);
HA h19_31(X31Y19,c18_31,c19_31,z19_31);
HA h20_31(X31Y20,c19_31,c20_31,z20_31);
HA h21_31(X31Y21,c20_31,c21_31,z21_31);
HA h22_31(X31Y22,c21_31,c22_31,z22_31);
HA h23_31(X31Y23,c22_31,c23_31,z23_31);
HA h24_31(X31Y24,c23_31,c24_31,z24_31);
HA h25_31(X31Y25,c24_31,c25_31,z25_31);
HA h26_31(X31Y26,c25_31,c26_31,z26_31);
HA h27_31(X31Y27,c26_31,c27_31,z27_31);
HA h28_31(X31Y28,c27_31,c28_31,z28_31);
HA h29_31(X31Y29,c28_31,c29_31,z29_31);
HA h30_31(X31Y30,c29_31,c30_31,z30_31);
HA h31_31(X31Y31,c30_31,c31_31,z31_31);
HA h32(z31_1,c31_0,c32,Z[32]);

assign z31_32 = 1;
FA f2_0(X0Y2,z1_1,c1_0,c2_0,z2_0);
FA f2_1(X1Y2,z1_2,c1_1,c2_1,z2_1);
FA f2_2(X2Y2,z1_3,c1_2,c2_2,z2_2);
FA f2_3(X3Y2,z1_4,c1_3,c2_3,z2_3);
FA f2_4(X4Y2,z1_5,c1_4,c2_4,z2_4);
FA f2_5(X5Y2,z1_6,c1_5,c2_5,z2_5);
FA f2_6(X6Y2,z1_7,c1_6,c2_6,z2_6);
FA f2_7(X7Y2,z1_8,c1_7,c2_7,z2_7);
FA f2_8(X8Y2,z1_9,c1_8,c2_8,z2_8);
FA f2_9(X9Y2,z1_10,c1_9,c2_9,z2_9);
FA f2_10(X10Y2,z1_11,c1_10,c2_10,z2_10);
FA f2_11(X11Y2,z1_12,c1_11,c2_11,z2_11);
FA f2_12(X12Y2,z1_13,c1_12,c2_12,z2_12);
FA f2_13(X13Y2,z1_14,c1_13,c2_13,z2_13);
FA f2_14(X14Y2,z1_15,c1_14,c2_14,z2_14);
FA f2_15(X15Y2,z1_16,c1_15,c2_15,z2_15);
FA f2_16(X16Y2,z1_17,c1_16,c2_16,z2_16);
FA f2_17(X17Y2,z1_18,c1_17,c2_17,z2_17);
FA f2_18(X18Y2,z1_19,c1_18,c2_18,z2_18);
FA f2_19(X19Y2,z1_20,c1_19,c2_19,z2_19);
FA f2_20(X20Y2,z1_21,c1_20,c2_20,z2_20);
FA f2_21(X21Y2,z1_22,c1_21,c2_21,z2_21);
FA f2_22(X22Y2,z1_23,c1_22,c2_22,z2_22);
FA f2_23(X23Y2,z1_24,c1_23,c2_23,z2_23);
FA f2_24(X24Y2,z1_25,c1_24,c2_24,z2_24);
FA f2_25(X25Y2,z1_26,c1_25,c2_25,z2_25);
FA f2_26(X26Y2,z1_27,c1_26,c2_26,z2_26);
FA f2_27(X27Y2,z1_28,c1_27,c2_27,z2_27);
FA f2_28(X28Y2,z1_29,c1_28,c2_28,z2_28);
FA f2_29(X29Y2,z1_30,c1_29,c2_29,z2_29);
FA f2_30(X30Y2,z1_31,c1_30,c2_30,z2_30);
FA f3_0(X0Y3,z2_1,c2_0,c3_0,z3_0);
FA f3_1(X1Y3,z2_2,c2_1,c3_1,z3_1);
FA f3_2(X2Y3,z2_3,c2_2,c3_2,z3_2);
FA f3_3(X3Y3,z2_4,c2_3,c3_3,z3_3);
FA f3_4(X4Y3,z2_5,c2_4,c3_4,z3_4);
FA f3_5(X5Y3,z2_6,c2_5,c3_5,z3_5);
FA f3_6(X6Y3,z2_7,c2_6,c3_6,z3_6);
FA f3_7(X7Y3,z2_8,c2_7,c3_7,z3_7);
FA f3_8(X8Y3,z2_9,c2_8,c3_8,z3_8);
FA f3_9(X9Y3,z2_10,c2_9,c3_9,z3_9);
FA f3_10(X10Y3,z2_11,c2_10,c3_10,z3_10);
FA f3_11(X11Y3,z2_12,c2_11,c3_11,z3_11);
FA f3_12(X12Y3,z2_13,c2_12,c3_12,z3_12);
FA f3_13(X13Y3,z2_14,c2_13,c3_13,z3_13);
FA f3_14(X14Y3,z2_15,c2_14,c3_14,z3_14);
FA f3_15(X15Y3,z2_16,c2_15,c3_15,z3_15);
FA f3_16(X16Y3,z2_17,c2_16,c3_16,z3_16);
FA f3_17(X17Y3,z2_18,c2_17,c3_17,z3_17);
FA f3_18(X18Y3,z2_19,c2_18,c3_18,z3_18);
FA f3_19(X19Y3,z2_20,c2_19,c3_19,z3_19);
FA f3_20(X20Y3,z2_21,c2_20,c3_20,z3_20);
FA f3_21(X21Y3,z2_22,c2_21,c3_21,z3_21);
FA f3_22(X22Y3,z2_23,c2_22,c3_22,z3_22);
FA f3_23(X23Y3,z2_24,c2_23,c3_23,z3_23);
FA f3_24(X24Y3,z2_25,c2_24,c3_24,z3_24);
FA f3_25(X25Y3,z2_26,c2_25,c3_25,z3_25);
FA f3_26(X26Y3,z2_27,c2_26,c3_26,z3_26);
FA f3_27(X27Y3,z2_28,c2_27,c3_27,z3_27);
FA f3_28(X28Y3,z2_29,c2_28,c3_28,z3_28);
FA f3_29(X29Y3,z2_30,c2_29,c3_29,z3_29);
FA f3_30(X30Y3,z2_31,c2_30,c3_30,z3_30);
FA f4_0(X0Y4,z3_1,c3_0,c4_0,z4_0);
FA f4_1(X1Y4,z3_2,c3_1,c4_1,z4_1);
FA f4_2(X2Y4,z3_3,c3_2,c4_2,z4_2);
FA f4_3(X3Y4,z3_4,c3_3,c4_3,z4_3);
FA f4_4(X4Y4,z3_5,c3_4,c4_4,z4_4);
FA f4_5(X5Y4,z3_6,c3_5,c4_5,z4_5);
FA f4_6(X6Y4,z3_7,c3_6,c4_6,z4_6);
FA f4_7(X7Y4,z3_8,c3_7,c4_7,z4_7);
FA f4_8(X8Y4,z3_9,c3_8,c4_8,z4_8);
FA f4_9(X9Y4,z3_10,c3_9,c4_9,z4_9);
FA f4_10(X10Y4,z3_11,c3_10,c4_10,z4_10);
FA f4_11(X11Y4,z3_12,c3_11,c4_11,z4_11);
FA f4_12(X12Y4,z3_13,c3_12,c4_12,z4_12);
FA f4_13(X13Y4,z3_14,c3_13,c4_13,z4_13);
FA f4_14(X14Y4,z3_15,c3_14,c4_14,z4_14);
FA f4_15(X15Y4,z3_16,c3_15,c4_15,z4_15);
FA f4_16(X16Y4,z3_17,c3_16,c4_16,z4_16);
FA f4_17(X17Y4,z3_18,c3_17,c4_17,z4_17);
FA f4_18(X18Y4,z3_19,c3_18,c4_18,z4_18);
FA f4_19(X19Y4,z3_20,c3_19,c4_19,z4_19);
FA f4_20(X20Y4,z3_21,c3_20,c4_20,z4_20);
FA f4_21(X21Y4,z3_22,c3_21,c4_21,z4_21);
FA f4_22(X22Y4,z3_23,c3_22,c4_22,z4_22);
FA f4_23(X23Y4,z3_24,c3_23,c4_23,z4_23);
FA f4_24(X24Y4,z3_25,c3_24,c4_24,z4_24);
FA f4_25(X25Y4,z3_26,c3_25,c4_25,z4_25);
FA f4_26(X26Y4,z3_27,c3_26,c4_26,z4_26);
FA f4_27(X27Y4,z3_28,c3_27,c4_27,z4_27);
FA f4_28(X28Y4,z3_29,c3_28,c4_28,z4_28);
FA f4_29(X29Y4,z3_30,c3_29,c4_29,z4_29);
FA f4_30(X30Y4,z3_31,c3_30,c4_30,z4_30);
FA f5_0(X0Y5,z4_1,c4_0,c5_0,z5_0);
FA f5_1(X1Y5,z4_2,c4_1,c5_1,z5_1);
FA f5_2(X2Y5,z4_3,c4_2,c5_2,z5_2);
FA f5_3(X3Y5,z4_4,c4_3,c5_3,z5_3);
FA f5_4(X4Y5,z4_5,c4_4,c5_4,z5_4);
FA f5_5(X5Y5,z4_6,c4_5,c5_5,z5_5);
FA f5_6(X6Y5,z4_7,c4_6,c5_6,z5_6);
FA f5_7(X7Y5,z4_8,c4_7,c5_7,z5_7);
FA f5_8(X8Y5,z4_9,c4_8,c5_8,z5_8);
FA f5_9(X9Y5,z4_10,c4_9,c5_9,z5_9);
FA f5_10(X10Y5,z4_11,c4_10,c5_10,z5_10);
FA f5_11(X11Y5,z4_12,c4_11,c5_11,z5_11);
FA f5_12(X12Y5,z4_13,c4_12,c5_12,z5_12);
FA f5_13(X13Y5,z4_14,c4_13,c5_13,z5_13);
FA f5_14(X14Y5,z4_15,c4_14,c5_14,z5_14);
FA f5_15(X15Y5,z4_16,c4_15,c5_15,z5_15);
FA f5_16(X16Y5,z4_17,c4_16,c5_16,z5_16);
FA f5_17(X17Y5,z4_18,c4_17,c5_17,z5_17);
FA f5_18(X18Y5,z4_19,c4_18,c5_18,z5_18);
FA f5_19(X19Y5,z4_20,c4_19,c5_19,z5_19);
FA f5_20(X20Y5,z4_21,c4_20,c5_20,z5_20);
FA f5_21(X21Y5,z4_22,c4_21,c5_21,z5_21);
FA f5_22(X22Y5,z4_23,c4_22,c5_22,z5_22);
FA f5_23(X23Y5,z4_24,c4_23,c5_23,z5_23);
FA f5_24(X24Y5,z4_25,c4_24,c5_24,z5_24);
FA f5_25(X25Y5,z4_26,c4_25,c5_25,z5_25);
FA f5_26(X26Y5,z4_27,c4_26,c5_26,z5_26);
FA f5_27(X27Y5,z4_28,c4_27,c5_27,z5_27);
FA f5_28(X28Y5,z4_29,c4_28,c5_28,z5_28);
FA f5_29(X29Y5,z4_30,c4_29,c5_29,z5_29);
FA f5_30(X30Y5,z4_31,c4_30,c5_30,z5_30);
FA f6_0(X0Y6,z5_1,c5_0,c6_0,z6_0);
FA f6_1(X1Y6,z5_2,c5_1,c6_1,z6_1);
FA f6_2(X2Y6,z5_3,c5_2,c6_2,z6_2);
FA f6_3(X3Y6,z5_4,c5_3,c6_3,z6_3);
FA f6_4(X4Y6,z5_5,c5_4,c6_4,z6_4);
FA f6_5(X5Y6,z5_6,c5_5,c6_5,z6_5);
FA f6_6(X6Y6,z5_7,c5_6,c6_6,z6_6);
FA f6_7(X7Y6,z5_8,c5_7,c6_7,z6_7);
FA f6_8(X8Y6,z5_9,c5_8,c6_8,z6_8);
FA f6_9(X9Y6,z5_10,c5_9,c6_9,z6_9);
FA f6_10(X10Y6,z5_11,c5_10,c6_10,z6_10);
FA f6_11(X11Y6,z5_12,c5_11,c6_11,z6_11);
FA f6_12(X12Y6,z5_13,c5_12,c6_12,z6_12);
FA f6_13(X13Y6,z5_14,c5_13,c6_13,z6_13);
FA f6_14(X14Y6,z5_15,c5_14,c6_14,z6_14);
FA f6_15(X15Y6,z5_16,c5_15,c6_15,z6_15);
FA f6_16(X16Y6,z5_17,c5_16,c6_16,z6_16);
FA f6_17(X17Y6,z5_18,c5_17,c6_17,z6_17);
FA f6_18(X18Y6,z5_19,c5_18,c6_18,z6_18);
FA f6_19(X19Y6,z5_20,c5_19,c6_19,z6_19);
FA f6_20(X20Y6,z5_21,c5_20,c6_20,z6_20);
FA f6_21(X21Y6,z5_22,c5_21,c6_21,z6_21);
FA f6_22(X22Y6,z5_23,c5_22,c6_22,z6_22);
FA f6_23(X23Y6,z5_24,c5_23,c6_23,z6_23);
FA f6_24(X24Y6,z5_25,c5_24,c6_24,z6_24);
FA f6_25(X25Y6,z5_26,c5_25,c6_25,z6_25);
FA f6_26(X26Y6,z5_27,c5_26,c6_26,z6_26);
FA f6_27(X27Y6,z5_28,c5_27,c6_27,z6_27);
FA f6_28(X28Y6,z5_29,c5_28,c6_28,z6_28);
FA f6_29(X29Y6,z5_30,c5_29,c6_29,z6_29);
FA f6_30(X30Y6,z5_31,c5_30,c6_30,z6_30);
FA f7_0(X0Y7,z6_1,c6_0,c7_0,z7_0);
FA f7_1(X1Y7,z6_2,c6_1,c7_1,z7_1);
FA f7_2(X2Y7,z6_3,c6_2,c7_2,z7_2);
FA f7_3(X3Y7,z6_4,c6_3,c7_3,z7_3);
FA f7_4(X4Y7,z6_5,c6_4,c7_4,z7_4);
FA f7_5(X5Y7,z6_6,c6_5,c7_5,z7_5);
FA f7_6(X6Y7,z6_7,c6_6,c7_6,z7_6);
FA f7_7(X7Y7,z6_8,c6_7,c7_7,z7_7);
FA f7_8(X8Y7,z6_9,c6_8,c7_8,z7_8);
FA f7_9(X9Y7,z6_10,c6_9,c7_9,z7_9);
FA f7_10(X10Y7,z6_11,c6_10,c7_10,z7_10);
FA f7_11(X11Y7,z6_12,c6_11,c7_11,z7_11);
FA f7_12(X12Y7,z6_13,c6_12,c7_12,z7_12);
FA f7_13(X13Y7,z6_14,c6_13,c7_13,z7_13);
FA f7_14(X14Y7,z6_15,c6_14,c7_14,z7_14);
FA f7_15(X15Y7,z6_16,c6_15,c7_15,z7_15);
FA f7_16(X16Y7,z6_17,c6_16,c7_16,z7_16);
FA f7_17(X17Y7,z6_18,c6_17,c7_17,z7_17);
FA f7_18(X18Y7,z6_19,c6_18,c7_18,z7_18);
FA f7_19(X19Y7,z6_20,c6_19,c7_19,z7_19);
FA f7_20(X20Y7,z6_21,c6_20,c7_20,z7_20);
FA f7_21(X21Y7,z6_22,c6_21,c7_21,z7_21);
FA f7_22(X22Y7,z6_23,c6_22,c7_22,z7_22);
FA f7_23(X23Y7,z6_24,c6_23,c7_23,z7_23);
FA f7_24(X24Y7,z6_25,c6_24,c7_24,z7_24);
FA f7_25(X25Y7,z6_26,c6_25,c7_25,z7_25);
FA f7_26(X26Y7,z6_27,c6_26,c7_26,z7_26);
FA f7_27(X27Y7,z6_28,c6_27,c7_27,z7_27);
FA f7_28(X28Y7,z6_29,c6_28,c7_28,z7_28);
FA f7_29(X29Y7,z6_30,c6_29,c7_29,z7_29);
FA f7_30(X30Y7,z6_31,c6_30,c7_30,z7_30);
FA f8_0(X0Y8,z7_1,c7_0,c8_0,z8_0);
FA f8_1(X1Y8,z7_2,c7_1,c8_1,z8_1);
FA f8_2(X2Y8,z7_3,c7_2,c8_2,z8_2);
FA f8_3(X3Y8,z7_4,c7_3,c8_3,z8_3);
FA f8_4(X4Y8,z7_5,c7_4,c8_4,z8_4);
FA f8_5(X5Y8,z7_6,c7_5,c8_5,z8_5);
FA f8_6(X6Y8,z7_7,c7_6,c8_6,z8_6);
FA f8_7(X7Y8,z7_8,c7_7,c8_7,z8_7);
FA f8_8(X8Y8,z7_9,c7_8,c8_8,z8_8);
FA f8_9(X9Y8,z7_10,c7_9,c8_9,z8_9);
FA f8_10(X10Y8,z7_11,c7_10,c8_10,z8_10);
FA f8_11(X11Y8,z7_12,c7_11,c8_11,z8_11);
FA f8_12(X12Y8,z7_13,c7_12,c8_12,z8_12);
FA f8_13(X13Y8,z7_14,c7_13,c8_13,z8_13);
FA f8_14(X14Y8,z7_15,c7_14,c8_14,z8_14);
FA f8_15(X15Y8,z7_16,c7_15,c8_15,z8_15);
FA f8_16(X16Y8,z7_17,c7_16,c8_16,z8_16);
FA f8_17(X17Y8,z7_18,c7_17,c8_17,z8_17);
FA f8_18(X18Y8,z7_19,c7_18,c8_18,z8_18);
FA f8_19(X19Y8,z7_20,c7_19,c8_19,z8_19);
FA f8_20(X20Y8,z7_21,c7_20,c8_20,z8_20);
FA f8_21(X21Y8,z7_22,c7_21,c8_21,z8_21);
FA f8_22(X22Y8,z7_23,c7_22,c8_22,z8_22);
FA f8_23(X23Y8,z7_24,c7_23,c8_23,z8_23);
FA f8_24(X24Y8,z7_25,c7_24,c8_24,z8_24);
FA f8_25(X25Y8,z7_26,c7_25,c8_25,z8_25);
FA f8_26(X26Y8,z7_27,c7_26,c8_26,z8_26);
FA f8_27(X27Y8,z7_28,c7_27,c8_27,z8_27);
FA f8_28(X28Y8,z7_29,c7_28,c8_28,z8_28);
FA f8_29(X29Y8,z7_30,c7_29,c8_29,z8_29);
FA f8_30(X30Y8,z7_31,c7_30,c8_30,z8_30);
FA f9_0(X0Y9,z8_1,c8_0,c9_0,z9_0);
FA f9_1(X1Y9,z8_2,c8_1,c9_1,z9_1);
FA f9_2(X2Y9,z8_3,c8_2,c9_2,z9_2);
FA f9_3(X3Y9,z8_4,c8_3,c9_3,z9_3);
FA f9_4(X4Y9,z8_5,c8_4,c9_4,z9_4);
FA f9_5(X5Y9,z8_6,c8_5,c9_5,z9_5);
FA f9_6(X6Y9,z8_7,c8_6,c9_6,z9_6);
FA f9_7(X7Y9,z8_8,c8_7,c9_7,z9_7);
FA f9_8(X8Y9,z8_9,c8_8,c9_8,z9_8);
FA f9_9(X9Y9,z8_10,c8_9,c9_9,z9_9);
FA f9_10(X10Y9,z8_11,c8_10,c9_10,z9_10);
FA f9_11(X11Y9,z8_12,c8_11,c9_11,z9_11);
FA f9_12(X12Y9,z8_13,c8_12,c9_12,z9_12);
FA f9_13(X13Y9,z8_14,c8_13,c9_13,z9_13);
FA f9_14(X14Y9,z8_15,c8_14,c9_14,z9_14);
FA f9_15(X15Y9,z8_16,c8_15,c9_15,z9_15);
FA f9_16(X16Y9,z8_17,c8_16,c9_16,z9_16);
FA f9_17(X17Y9,z8_18,c8_17,c9_17,z9_17);
FA f9_18(X18Y9,z8_19,c8_18,c9_18,z9_18);
FA f9_19(X19Y9,z8_20,c8_19,c9_19,z9_19);
FA f9_20(X20Y9,z8_21,c8_20,c9_20,z9_20);
FA f9_21(X21Y9,z8_22,c8_21,c9_21,z9_21);
FA f9_22(X22Y9,z8_23,c8_22,c9_22,z9_22);
FA f9_23(X23Y9,z8_24,c8_23,c9_23,z9_23);
FA f9_24(X24Y9,z8_25,c8_24,c9_24,z9_24);
FA f9_25(X25Y9,z8_26,c8_25,c9_25,z9_25);
FA f9_26(X26Y9,z8_27,c8_26,c9_26,z9_26);
FA f9_27(X27Y9,z8_28,c8_27,c9_27,z9_27);
FA f9_28(X28Y9,z8_29,c8_28,c9_28,z9_28);
FA f9_29(X29Y9,z8_30,c8_29,c9_29,z9_29);
FA f9_30(X30Y9,z8_31,c8_30,c9_30,z9_30);
FA f10_0(X0Y10,z9_1,c9_0,c10_0,z10_0);
FA f10_1(X1Y10,z9_2,c9_1,c10_1,z10_1);
FA f10_2(X2Y10,z9_3,c9_2,c10_2,z10_2);
FA f10_3(X3Y10,z9_4,c9_3,c10_3,z10_3);
FA f10_4(X4Y10,z9_5,c9_4,c10_4,z10_4);
FA f10_5(X5Y10,z9_6,c9_5,c10_5,z10_5);
FA f10_6(X6Y10,z9_7,c9_6,c10_6,z10_6);
FA f10_7(X7Y10,z9_8,c9_7,c10_7,z10_7);
FA f10_8(X8Y10,z9_9,c9_8,c10_8,z10_8);
FA f10_9(X9Y10,z9_10,c9_9,c10_9,z10_9);
FA f10_10(X10Y10,z9_11,c9_10,c10_10,z10_10);
FA f10_11(X11Y10,z9_12,c9_11,c10_11,z10_11);
FA f10_12(X12Y10,z9_13,c9_12,c10_12,z10_12);
FA f10_13(X13Y10,z9_14,c9_13,c10_13,z10_13);
FA f10_14(X14Y10,z9_15,c9_14,c10_14,z10_14);
FA f10_15(X15Y10,z9_16,c9_15,c10_15,z10_15);
FA f10_16(X16Y10,z9_17,c9_16,c10_16,z10_16);
FA f10_17(X17Y10,z9_18,c9_17,c10_17,z10_17);
FA f10_18(X18Y10,z9_19,c9_18,c10_18,z10_18);
FA f10_19(X19Y10,z9_20,c9_19,c10_19,z10_19);
FA f10_20(X20Y10,z9_21,c9_20,c10_20,z10_20);
FA f10_21(X21Y10,z9_22,c9_21,c10_21,z10_21);
FA f10_22(X22Y10,z9_23,c9_22,c10_22,z10_22);
FA f10_23(X23Y10,z9_24,c9_23,c10_23,z10_23);
FA f10_24(X24Y10,z9_25,c9_24,c10_24,z10_24);
FA f10_25(X25Y10,z9_26,c9_25,c10_25,z10_25);
FA f10_26(X26Y10,z9_27,c9_26,c10_26,z10_26);
FA f10_27(X27Y10,z9_28,c9_27,c10_27,z10_27);
FA f10_28(X28Y10,z9_29,c9_28,c10_28,z10_28);
FA f10_29(X29Y10,z9_30,c9_29,c10_29,z10_29);
FA f10_30(X30Y10,z9_31,c9_30,c10_30,z10_30);
FA f11_0(X0Y11,z10_1,c10_0,c11_0,z11_0);
FA f11_1(X1Y11,z10_2,c10_1,c11_1,z11_1);
FA f11_2(X2Y11,z10_3,c10_2,c11_2,z11_2);
FA f11_3(X3Y11,z10_4,c10_3,c11_3,z11_3);
FA f11_4(X4Y11,z10_5,c10_4,c11_4,z11_4);
FA f11_5(X5Y11,z10_6,c10_5,c11_5,z11_5);
FA f11_6(X6Y11,z10_7,c10_6,c11_6,z11_6);
FA f11_7(X7Y11,z10_8,c10_7,c11_7,z11_7);
FA f11_8(X8Y11,z10_9,c10_8,c11_8,z11_8);
FA f11_9(X9Y11,z10_10,c10_9,c11_9,z11_9);
FA f11_10(X10Y11,z10_11,c10_10,c11_10,z11_10);
FA f11_11(X11Y11,z10_12,c10_11,c11_11,z11_11);
FA f11_12(X12Y11,z10_13,c10_12,c11_12,z11_12);
FA f11_13(X13Y11,z10_14,c10_13,c11_13,z11_13);
FA f11_14(X14Y11,z10_15,c10_14,c11_14,z11_14);
FA f11_15(X15Y11,z10_16,c10_15,c11_15,z11_15);
FA f11_16(X16Y11,z10_17,c10_16,c11_16,z11_16);
FA f11_17(X17Y11,z10_18,c10_17,c11_17,z11_17);
FA f11_18(X18Y11,z10_19,c10_18,c11_18,z11_18);
FA f11_19(X19Y11,z10_20,c10_19,c11_19,z11_19);
FA f11_20(X20Y11,z10_21,c10_20,c11_20,z11_20);
FA f11_21(X21Y11,z10_22,c10_21,c11_21,z11_21);
FA f11_22(X22Y11,z10_23,c10_22,c11_22,z11_22);
FA f11_23(X23Y11,z10_24,c10_23,c11_23,z11_23);
FA f11_24(X24Y11,z10_25,c10_24,c11_24,z11_24);
FA f11_25(X25Y11,z10_26,c10_25,c11_25,z11_25);
FA f11_26(X26Y11,z10_27,c10_26,c11_26,z11_26);
FA f11_27(X27Y11,z10_28,c10_27,c11_27,z11_27);
FA f11_28(X28Y11,z10_29,c10_28,c11_28,z11_28);
FA f11_29(X29Y11,z10_30,c10_29,c11_29,z11_29);
FA f11_30(X30Y11,z10_31,c10_30,c11_30,z11_30);
FA f12_0(X0Y12,z11_1,c11_0,c12_0,z12_0);
FA f12_1(X1Y12,z11_2,c11_1,c12_1,z12_1);
FA f12_2(X2Y12,z11_3,c11_2,c12_2,z12_2);
FA f12_3(X3Y12,z11_4,c11_3,c12_3,z12_3);
FA f12_4(X4Y12,z11_5,c11_4,c12_4,z12_4);
FA f12_5(X5Y12,z11_6,c11_5,c12_5,z12_5);
FA f12_6(X6Y12,z11_7,c11_6,c12_6,z12_6);
FA f12_7(X7Y12,z11_8,c11_7,c12_7,z12_7);
FA f12_8(X8Y12,z11_9,c11_8,c12_8,z12_8);
FA f12_9(X9Y12,z11_10,c11_9,c12_9,z12_9);
FA f12_10(X10Y12,z11_11,c11_10,c12_10,z12_10);
FA f12_11(X11Y12,z11_12,c11_11,c12_11,z12_11);
FA f12_12(X12Y12,z11_13,c11_12,c12_12,z12_12);
FA f12_13(X13Y12,z11_14,c11_13,c12_13,z12_13);
FA f12_14(X14Y12,z11_15,c11_14,c12_14,z12_14);
FA f12_15(X15Y12,z11_16,c11_15,c12_15,z12_15);
FA f12_16(X16Y12,z11_17,c11_16,c12_16,z12_16);
FA f12_17(X17Y12,z11_18,c11_17,c12_17,z12_17);
FA f12_18(X18Y12,z11_19,c11_18,c12_18,z12_18);
FA f12_19(X19Y12,z11_20,c11_19,c12_19,z12_19);
FA f12_20(X20Y12,z11_21,c11_20,c12_20,z12_20);
FA f12_21(X21Y12,z11_22,c11_21,c12_21,z12_21);
FA f12_22(X22Y12,z11_23,c11_22,c12_22,z12_22);
FA f12_23(X23Y12,z11_24,c11_23,c12_23,z12_23);
FA f12_24(X24Y12,z11_25,c11_24,c12_24,z12_24);
FA f12_25(X25Y12,z11_26,c11_25,c12_25,z12_25);
FA f12_26(X26Y12,z11_27,c11_26,c12_26,z12_26);
FA f12_27(X27Y12,z11_28,c11_27,c12_27,z12_27);
FA f12_28(X28Y12,z11_29,c11_28,c12_28,z12_28);
FA f12_29(X29Y12,z11_30,c11_29,c12_29,z12_29);
FA f12_30(X30Y12,z11_31,c11_30,c12_30,z12_30);
FA f13_0(X0Y13,z12_1,c12_0,c13_0,z13_0);
FA f13_1(X1Y13,z12_2,c12_1,c13_1,z13_1);
FA f13_2(X2Y13,z12_3,c12_2,c13_2,z13_2);
FA f13_3(X3Y13,z12_4,c12_3,c13_3,z13_3);
FA f13_4(X4Y13,z12_5,c12_4,c13_4,z13_4);
FA f13_5(X5Y13,z12_6,c12_5,c13_5,z13_5);
FA f13_6(X6Y13,z12_7,c12_6,c13_6,z13_6);
FA f13_7(X7Y13,z12_8,c12_7,c13_7,z13_7);
FA f13_8(X8Y13,z12_9,c12_8,c13_8,z13_8);
FA f13_9(X9Y13,z12_10,c12_9,c13_9,z13_9);
FA f13_10(X10Y13,z12_11,c12_10,c13_10,z13_10);
FA f13_11(X11Y13,z12_12,c12_11,c13_11,z13_11);
FA f13_12(X12Y13,z12_13,c12_12,c13_12,z13_12);
FA f13_13(X13Y13,z12_14,c12_13,c13_13,z13_13);
FA f13_14(X14Y13,z12_15,c12_14,c13_14,z13_14);
FA f13_15(X15Y13,z12_16,c12_15,c13_15,z13_15);
FA f13_16(X16Y13,z12_17,c12_16,c13_16,z13_16);
FA f13_17(X17Y13,z12_18,c12_17,c13_17,z13_17);
FA f13_18(X18Y13,z12_19,c12_18,c13_18,z13_18);
FA f13_19(X19Y13,z12_20,c12_19,c13_19,z13_19);
FA f13_20(X20Y13,z12_21,c12_20,c13_20,z13_20);
FA f13_21(X21Y13,z12_22,c12_21,c13_21,z13_21);
FA f13_22(X22Y13,z12_23,c12_22,c13_22,z13_22);
FA f13_23(X23Y13,z12_24,c12_23,c13_23,z13_23);
FA f13_24(X24Y13,z12_25,c12_24,c13_24,z13_24);
FA f13_25(X25Y13,z12_26,c12_25,c13_25,z13_25);
FA f13_26(X26Y13,z12_27,c12_26,c13_26,z13_26);
FA f13_27(X27Y13,z12_28,c12_27,c13_27,z13_27);
FA f13_28(X28Y13,z12_29,c12_28,c13_28,z13_28);
FA f13_29(X29Y13,z12_30,c12_29,c13_29,z13_29);
FA f13_30(X30Y13,z12_31,c12_30,c13_30,z13_30);
FA f14_0(X0Y14,z13_1,c13_0,c14_0,z14_0);
FA f14_1(X1Y14,z13_2,c13_1,c14_1,z14_1);
FA f14_2(X2Y14,z13_3,c13_2,c14_2,z14_2);
FA f14_3(X3Y14,z13_4,c13_3,c14_3,z14_3);
FA f14_4(X4Y14,z13_5,c13_4,c14_4,z14_4);
FA f14_5(X5Y14,z13_6,c13_5,c14_5,z14_5);
FA f14_6(X6Y14,z13_7,c13_6,c14_6,z14_6);
FA f14_7(X7Y14,z13_8,c13_7,c14_7,z14_7);
FA f14_8(X8Y14,z13_9,c13_8,c14_8,z14_8);
FA f14_9(X9Y14,z13_10,c13_9,c14_9,z14_9);
FA f14_10(X10Y14,z13_11,c13_10,c14_10,z14_10);
FA f14_11(X11Y14,z13_12,c13_11,c14_11,z14_11);
FA f14_12(X12Y14,z13_13,c13_12,c14_12,z14_12);
FA f14_13(X13Y14,z13_14,c13_13,c14_13,z14_13);
FA f14_14(X14Y14,z13_15,c13_14,c14_14,z14_14);
FA f14_15(X15Y14,z13_16,c13_15,c14_15,z14_15);
FA f14_16(X16Y14,z13_17,c13_16,c14_16,z14_16);
FA f14_17(X17Y14,z13_18,c13_17,c14_17,z14_17);
FA f14_18(X18Y14,z13_19,c13_18,c14_18,z14_18);
FA f14_19(X19Y14,z13_20,c13_19,c14_19,z14_19);
FA f14_20(X20Y14,z13_21,c13_20,c14_20,z14_20);
FA f14_21(X21Y14,z13_22,c13_21,c14_21,z14_21);
FA f14_22(X22Y14,z13_23,c13_22,c14_22,z14_22);
FA f14_23(X23Y14,z13_24,c13_23,c14_23,z14_23);
FA f14_24(X24Y14,z13_25,c13_24,c14_24,z14_24);
FA f14_25(X25Y14,z13_26,c13_25,c14_25,z14_25);
FA f14_26(X26Y14,z13_27,c13_26,c14_26,z14_26);
FA f14_27(X27Y14,z13_28,c13_27,c14_27,z14_27);
FA f14_28(X28Y14,z13_29,c13_28,c14_28,z14_28);
FA f14_29(X29Y14,z13_30,c13_29,c14_29,z14_29);
FA f14_30(X30Y14,z13_31,c13_30,c14_30,z14_30);
FA f15_0(X0Y15,z14_1,c14_0,c15_0,z15_0);
FA f15_1(X1Y15,z14_2,c14_1,c15_1,z15_1);
FA f15_2(X2Y15,z14_3,c14_2,c15_2,z15_2);
FA f15_3(X3Y15,z14_4,c14_3,c15_3,z15_3);
FA f15_4(X4Y15,z14_5,c14_4,c15_4,z15_4);
FA f15_5(X5Y15,z14_6,c14_5,c15_5,z15_5);
FA f15_6(X6Y15,z14_7,c14_6,c15_6,z15_6);
FA f15_7(X7Y15,z14_8,c14_7,c15_7,z15_7);
FA f15_8(X8Y15,z14_9,c14_8,c15_8,z15_8);
FA f15_9(X9Y15,z14_10,c14_9,c15_9,z15_9);
FA f15_10(X10Y15,z14_11,c14_10,c15_10,z15_10);
FA f15_11(X11Y15,z14_12,c14_11,c15_11,z15_11);
FA f15_12(X12Y15,z14_13,c14_12,c15_12,z15_12);
FA f15_13(X13Y15,z14_14,c14_13,c15_13,z15_13);
FA f15_14(X14Y15,z14_15,c14_14,c15_14,z15_14);
FA f15_15(X15Y15,z14_16,c14_15,c15_15,z15_15);
FA f15_16(X16Y15,z14_17,c14_16,c15_16,z15_16);
FA f15_17(X17Y15,z14_18,c14_17,c15_17,z15_17);
FA f15_18(X18Y15,z14_19,c14_18,c15_18,z15_18);
FA f15_19(X19Y15,z14_20,c14_19,c15_19,z15_19);
FA f15_20(X20Y15,z14_21,c14_20,c15_20,z15_20);
FA f15_21(X21Y15,z14_22,c14_21,c15_21,z15_21);
FA f15_22(X22Y15,z14_23,c14_22,c15_22,z15_22);
FA f15_23(X23Y15,z14_24,c14_23,c15_23,z15_23);
FA f15_24(X24Y15,z14_25,c14_24,c15_24,z15_24);
FA f15_25(X25Y15,z14_26,c14_25,c15_25,z15_25);
FA f15_26(X26Y15,z14_27,c14_26,c15_26,z15_26);
FA f15_27(X27Y15,z14_28,c14_27,c15_27,z15_27);
FA f15_28(X28Y15,z14_29,c14_28,c15_28,z15_28);
FA f15_29(X29Y15,z14_30,c14_29,c15_29,z15_29);
FA f15_30(X30Y15,z14_31,c14_30,c15_30,z15_30);
FA f16_0(X0Y16,z15_1,c15_0,c16_0,z16_0);
FA f16_1(X1Y16,z15_2,c15_1,c16_1,z16_1);
FA f16_2(X2Y16,z15_3,c15_2,c16_2,z16_2);
FA f16_3(X3Y16,z15_4,c15_3,c16_3,z16_3);
FA f16_4(X4Y16,z15_5,c15_4,c16_4,z16_4);
FA f16_5(X5Y16,z15_6,c15_5,c16_5,z16_5);
FA f16_6(X6Y16,z15_7,c15_6,c16_6,z16_6);
FA f16_7(X7Y16,z15_8,c15_7,c16_7,z16_7);
FA f16_8(X8Y16,z15_9,c15_8,c16_8,z16_8);
FA f16_9(X9Y16,z15_10,c15_9,c16_9,z16_9);
FA f16_10(X10Y16,z15_11,c15_10,c16_10,z16_10);
FA f16_11(X11Y16,z15_12,c15_11,c16_11,z16_11);
FA f16_12(X12Y16,z15_13,c15_12,c16_12,z16_12);
FA f16_13(X13Y16,z15_14,c15_13,c16_13,z16_13);
FA f16_14(X14Y16,z15_15,c15_14,c16_14,z16_14);
FA f16_15(X15Y16,z15_16,c15_15,c16_15,z16_15);
FA f16_16(X16Y16,z15_17,c15_16,c16_16,z16_16);
FA f16_17(X17Y16,z15_18,c15_17,c16_17,z16_17);
FA f16_18(X18Y16,z15_19,c15_18,c16_18,z16_18);
FA f16_19(X19Y16,z15_20,c15_19,c16_19,z16_19);
FA f16_20(X20Y16,z15_21,c15_20,c16_20,z16_20);
FA f16_21(X21Y16,z15_22,c15_21,c16_21,z16_21);
FA f16_22(X22Y16,z15_23,c15_22,c16_22,z16_22);
FA f16_23(X23Y16,z15_24,c15_23,c16_23,z16_23);
FA f16_24(X24Y16,z15_25,c15_24,c16_24,z16_24);
FA f16_25(X25Y16,z15_26,c15_25,c16_25,z16_25);
FA f16_26(X26Y16,z15_27,c15_26,c16_26,z16_26);
FA f16_27(X27Y16,z15_28,c15_27,c16_27,z16_27);
FA f16_28(X28Y16,z15_29,c15_28,c16_28,z16_28);
FA f16_29(X29Y16,z15_30,c15_29,c16_29,z16_29);
FA f16_30(X30Y16,z15_31,c15_30,c16_30,z16_30);
FA f17_0(X0Y17,z16_1,c16_0,c17_0,z17_0);
FA f17_1(X1Y17,z16_2,c16_1,c17_1,z17_1);
FA f17_2(X2Y17,z16_3,c16_2,c17_2,z17_2);
FA f17_3(X3Y17,z16_4,c16_3,c17_3,z17_3);
FA f17_4(X4Y17,z16_5,c16_4,c17_4,z17_4);
FA f17_5(X5Y17,z16_6,c16_5,c17_5,z17_5);
FA f17_6(X6Y17,z16_7,c16_6,c17_6,z17_6);
FA f17_7(X7Y17,z16_8,c16_7,c17_7,z17_7);
FA f17_8(X8Y17,z16_9,c16_8,c17_8,z17_8);
FA f17_9(X9Y17,z16_10,c16_9,c17_9,z17_9);
FA f17_10(X10Y17,z16_11,c16_10,c17_10,z17_10);
FA f17_11(X11Y17,z16_12,c16_11,c17_11,z17_11);
FA f17_12(X12Y17,z16_13,c16_12,c17_12,z17_12);
FA f17_13(X13Y17,z16_14,c16_13,c17_13,z17_13);
FA f17_14(X14Y17,z16_15,c16_14,c17_14,z17_14);
FA f17_15(X15Y17,z16_16,c16_15,c17_15,z17_15);
FA f17_16(X16Y17,z16_17,c16_16,c17_16,z17_16);
FA f17_17(X17Y17,z16_18,c16_17,c17_17,z17_17);
FA f17_18(X18Y17,z16_19,c16_18,c17_18,z17_18);
FA f17_19(X19Y17,z16_20,c16_19,c17_19,z17_19);
FA f17_20(X20Y17,z16_21,c16_20,c17_20,z17_20);
FA f17_21(X21Y17,z16_22,c16_21,c17_21,z17_21);
FA f17_22(X22Y17,z16_23,c16_22,c17_22,z17_22);
FA f17_23(X23Y17,z16_24,c16_23,c17_23,z17_23);
FA f17_24(X24Y17,z16_25,c16_24,c17_24,z17_24);
FA f17_25(X25Y17,z16_26,c16_25,c17_25,z17_25);
FA f17_26(X26Y17,z16_27,c16_26,c17_26,z17_26);
FA f17_27(X27Y17,z16_28,c16_27,c17_27,z17_27);
FA f17_28(X28Y17,z16_29,c16_28,c17_28,z17_28);
FA f17_29(X29Y17,z16_30,c16_29,c17_29,z17_29);
FA f17_30(X30Y17,z16_31,c16_30,c17_30,z17_30);
FA f18_0(X0Y18,z17_1,c17_0,c18_0,z18_0);
FA f18_1(X1Y18,z17_2,c17_1,c18_1,z18_1);
FA f18_2(X2Y18,z17_3,c17_2,c18_2,z18_2);
FA f18_3(X3Y18,z17_4,c17_3,c18_3,z18_3);
FA f18_4(X4Y18,z17_5,c17_4,c18_4,z18_4);
FA f18_5(X5Y18,z17_6,c17_5,c18_5,z18_5);
FA f18_6(X6Y18,z17_7,c17_6,c18_6,z18_6);
FA f18_7(X7Y18,z17_8,c17_7,c18_7,z18_7);
FA f18_8(X8Y18,z17_9,c17_8,c18_8,z18_8);
FA f18_9(X9Y18,z17_10,c17_9,c18_9,z18_9);
FA f18_10(X10Y18,z17_11,c17_10,c18_10,z18_10);
FA f18_11(X11Y18,z17_12,c17_11,c18_11,z18_11);
FA f18_12(X12Y18,z17_13,c17_12,c18_12,z18_12);
FA f18_13(X13Y18,z17_14,c17_13,c18_13,z18_13);
FA f18_14(X14Y18,z17_15,c17_14,c18_14,z18_14);
FA f18_15(X15Y18,z17_16,c17_15,c18_15,z18_15);
FA f18_16(X16Y18,z17_17,c17_16,c18_16,z18_16);
FA f18_17(X17Y18,z17_18,c17_17,c18_17,z18_17);
FA f18_18(X18Y18,z17_19,c17_18,c18_18,z18_18);
FA f18_19(X19Y18,z17_20,c17_19,c18_19,z18_19);
FA f18_20(X20Y18,z17_21,c17_20,c18_20,z18_20);
FA f18_21(X21Y18,z17_22,c17_21,c18_21,z18_21);
FA f18_22(X22Y18,z17_23,c17_22,c18_22,z18_22);
FA f18_23(X23Y18,z17_24,c17_23,c18_23,z18_23);
FA f18_24(X24Y18,z17_25,c17_24,c18_24,z18_24);
FA f18_25(X25Y18,z17_26,c17_25,c18_25,z18_25);
FA f18_26(X26Y18,z17_27,c17_26,c18_26,z18_26);
FA f18_27(X27Y18,z17_28,c17_27,c18_27,z18_27);
FA f18_28(X28Y18,z17_29,c17_28,c18_28,z18_28);
FA f18_29(X29Y18,z17_30,c17_29,c18_29,z18_29);
FA f18_30(X30Y18,z17_31,c17_30,c18_30,z18_30);
FA f19_0(X0Y19,z18_1,c18_0,c19_0,z19_0);
FA f19_1(X1Y19,z18_2,c18_1,c19_1,z19_1);
FA f19_2(X2Y19,z18_3,c18_2,c19_2,z19_2);
FA f19_3(X3Y19,z18_4,c18_3,c19_3,z19_3);
FA f19_4(X4Y19,z18_5,c18_4,c19_4,z19_4);
FA f19_5(X5Y19,z18_6,c18_5,c19_5,z19_5);
FA f19_6(X6Y19,z18_7,c18_6,c19_6,z19_6);
FA f19_7(X7Y19,z18_8,c18_7,c19_7,z19_7);
FA f19_8(X8Y19,z18_9,c18_8,c19_8,z19_8);
FA f19_9(X9Y19,z18_10,c18_9,c19_9,z19_9);
FA f19_10(X10Y19,z18_11,c18_10,c19_10,z19_10);
FA f19_11(X11Y19,z18_12,c18_11,c19_11,z19_11);
FA f19_12(X12Y19,z18_13,c18_12,c19_12,z19_12);
FA f19_13(X13Y19,z18_14,c18_13,c19_13,z19_13);
FA f19_14(X14Y19,z18_15,c18_14,c19_14,z19_14);
FA f19_15(X15Y19,z18_16,c18_15,c19_15,z19_15);
FA f19_16(X16Y19,z18_17,c18_16,c19_16,z19_16);
FA f19_17(X17Y19,z18_18,c18_17,c19_17,z19_17);
FA f19_18(X18Y19,z18_19,c18_18,c19_18,z19_18);
FA f19_19(X19Y19,z18_20,c18_19,c19_19,z19_19);
FA f19_20(X20Y19,z18_21,c18_20,c19_20,z19_20);
FA f19_21(X21Y19,z18_22,c18_21,c19_21,z19_21);
FA f19_22(X22Y19,z18_23,c18_22,c19_22,z19_22);
FA f19_23(X23Y19,z18_24,c18_23,c19_23,z19_23);
FA f19_24(X24Y19,z18_25,c18_24,c19_24,z19_24);
FA f19_25(X25Y19,z18_26,c18_25,c19_25,z19_25);
FA f19_26(X26Y19,z18_27,c18_26,c19_26,z19_26);
FA f19_27(X27Y19,z18_28,c18_27,c19_27,z19_27);
FA f19_28(X28Y19,z18_29,c18_28,c19_28,z19_28);
FA f19_29(X29Y19,z18_30,c18_29,c19_29,z19_29);
FA f19_30(X30Y19,z18_31,c18_30,c19_30,z19_30);
FA f20_0(X0Y20,z19_1,c19_0,c20_0,z20_0);
FA f20_1(X1Y20,z19_2,c19_1,c20_1,z20_1);
FA f20_2(X2Y20,z19_3,c19_2,c20_2,z20_2);
FA f20_3(X3Y20,z19_4,c19_3,c20_3,z20_3);
FA f20_4(X4Y20,z19_5,c19_4,c20_4,z20_4);
FA f20_5(X5Y20,z19_6,c19_5,c20_5,z20_5);
FA f20_6(X6Y20,z19_7,c19_6,c20_6,z20_6);
FA f20_7(X7Y20,z19_8,c19_7,c20_7,z20_7);
FA f20_8(X8Y20,z19_9,c19_8,c20_8,z20_8);
FA f20_9(X9Y20,z19_10,c19_9,c20_9,z20_9);
FA f20_10(X10Y20,z19_11,c19_10,c20_10,z20_10);
FA f20_11(X11Y20,z19_12,c19_11,c20_11,z20_11);
FA f20_12(X12Y20,z19_13,c19_12,c20_12,z20_12);
FA f20_13(X13Y20,z19_14,c19_13,c20_13,z20_13);
FA f20_14(X14Y20,z19_15,c19_14,c20_14,z20_14);
FA f20_15(X15Y20,z19_16,c19_15,c20_15,z20_15);
FA f20_16(X16Y20,z19_17,c19_16,c20_16,z20_16);
FA f20_17(X17Y20,z19_18,c19_17,c20_17,z20_17);
FA f20_18(X18Y20,z19_19,c19_18,c20_18,z20_18);
FA f20_19(X19Y20,z19_20,c19_19,c20_19,z20_19);
FA f20_20(X20Y20,z19_21,c19_20,c20_20,z20_20);
FA f20_21(X21Y20,z19_22,c19_21,c20_21,z20_21);
FA f20_22(X22Y20,z19_23,c19_22,c20_22,z20_22);
FA f20_23(X23Y20,z19_24,c19_23,c20_23,z20_23);
FA f20_24(X24Y20,z19_25,c19_24,c20_24,z20_24);
FA f20_25(X25Y20,z19_26,c19_25,c20_25,z20_25);
FA f20_26(X26Y20,z19_27,c19_26,c20_26,z20_26);
FA f20_27(X27Y20,z19_28,c19_27,c20_27,z20_27);
FA f20_28(X28Y20,z19_29,c19_28,c20_28,z20_28);
FA f20_29(X29Y20,z19_30,c19_29,c20_29,z20_29);
FA f20_30(X30Y20,z19_31,c19_30,c20_30,z20_30);
FA f21_0(X0Y21,z20_1,c20_0,c21_0,z21_0);
FA f21_1(X1Y21,z20_2,c20_1,c21_1,z21_1);
FA f21_2(X2Y21,z20_3,c20_2,c21_2,z21_2);
FA f21_3(X3Y21,z20_4,c20_3,c21_3,z21_3);
FA f21_4(X4Y21,z20_5,c20_4,c21_4,z21_4);
FA f21_5(X5Y21,z20_6,c20_5,c21_5,z21_5);
FA f21_6(X6Y21,z20_7,c20_6,c21_6,z21_6);
FA f21_7(X7Y21,z20_8,c20_7,c21_7,z21_7);
FA f21_8(X8Y21,z20_9,c20_8,c21_8,z21_8);
FA f21_9(X9Y21,z20_10,c20_9,c21_9,z21_9);
FA f21_10(X10Y21,z20_11,c20_10,c21_10,z21_10);
FA f21_11(X11Y21,z20_12,c20_11,c21_11,z21_11);
FA f21_12(X12Y21,z20_13,c20_12,c21_12,z21_12);
FA f21_13(X13Y21,z20_14,c20_13,c21_13,z21_13);
FA f21_14(X14Y21,z20_15,c20_14,c21_14,z21_14);
FA f21_15(X15Y21,z20_16,c20_15,c21_15,z21_15);
FA f21_16(X16Y21,z20_17,c20_16,c21_16,z21_16);
FA f21_17(X17Y21,z20_18,c20_17,c21_17,z21_17);
FA f21_18(X18Y21,z20_19,c20_18,c21_18,z21_18);
FA f21_19(X19Y21,z20_20,c20_19,c21_19,z21_19);
FA f21_20(X20Y21,z20_21,c20_20,c21_20,z21_20);
FA f21_21(X21Y21,z20_22,c20_21,c21_21,z21_21);
FA f21_22(X22Y21,z20_23,c20_22,c21_22,z21_22);
FA f21_23(X23Y21,z20_24,c20_23,c21_23,z21_23);
FA f21_24(X24Y21,z20_25,c20_24,c21_24,z21_24);
FA f21_25(X25Y21,z20_26,c20_25,c21_25,z21_25);
FA f21_26(X26Y21,z20_27,c20_26,c21_26,z21_26);
FA f21_27(X27Y21,z20_28,c20_27,c21_27,z21_27);
FA f21_28(X28Y21,z20_29,c20_28,c21_28,z21_28);
FA f21_29(X29Y21,z20_30,c20_29,c21_29,z21_29);
FA f21_30(X30Y21,z20_31,c20_30,c21_30,z21_30);
FA f22_0(X0Y22,z21_1,c21_0,c22_0,z22_0);
FA f22_1(X1Y22,z21_2,c21_1,c22_1,z22_1);
FA f22_2(X2Y22,z21_3,c21_2,c22_2,z22_2);
FA f22_3(X3Y22,z21_4,c21_3,c22_3,z22_3);
FA f22_4(X4Y22,z21_5,c21_4,c22_4,z22_4);
FA f22_5(X5Y22,z21_6,c21_5,c22_5,z22_5);
FA f22_6(X6Y22,z21_7,c21_6,c22_6,z22_6);
FA f22_7(X7Y22,z21_8,c21_7,c22_7,z22_7);
FA f22_8(X8Y22,z21_9,c21_8,c22_8,z22_8);
FA f22_9(X9Y22,z21_10,c21_9,c22_9,z22_9);
FA f22_10(X10Y22,z21_11,c21_10,c22_10,z22_10);
FA f22_11(X11Y22,z21_12,c21_11,c22_11,z22_11);
FA f22_12(X12Y22,z21_13,c21_12,c22_12,z22_12);
FA f22_13(X13Y22,z21_14,c21_13,c22_13,z22_13);
FA f22_14(X14Y22,z21_15,c21_14,c22_14,z22_14);
FA f22_15(X15Y22,z21_16,c21_15,c22_15,z22_15);
FA f22_16(X16Y22,z21_17,c21_16,c22_16,z22_16);
FA f22_17(X17Y22,z21_18,c21_17,c22_17,z22_17);
FA f22_18(X18Y22,z21_19,c21_18,c22_18,z22_18);
FA f22_19(X19Y22,z21_20,c21_19,c22_19,z22_19);
FA f22_20(X20Y22,z21_21,c21_20,c22_20,z22_20);
FA f22_21(X21Y22,z21_22,c21_21,c22_21,z22_21);
FA f22_22(X22Y22,z21_23,c21_22,c22_22,z22_22);
FA f22_23(X23Y22,z21_24,c21_23,c22_23,z22_23);
FA f22_24(X24Y22,z21_25,c21_24,c22_24,z22_24);
FA f22_25(X25Y22,z21_26,c21_25,c22_25,z22_25);
FA f22_26(X26Y22,z21_27,c21_26,c22_26,z22_26);
FA f22_27(X27Y22,z21_28,c21_27,c22_27,z22_27);
FA f22_28(X28Y22,z21_29,c21_28,c22_28,z22_28);
FA f22_29(X29Y22,z21_30,c21_29,c22_29,z22_29);
FA f22_30(X30Y22,z21_31,c21_30,c22_30,z22_30);
FA f23_0(X0Y23,z22_1,c22_0,c23_0,z23_0);
FA f23_1(X1Y23,z22_2,c22_1,c23_1,z23_1);
FA f23_2(X2Y23,z22_3,c22_2,c23_2,z23_2);
FA f23_3(X3Y23,z22_4,c22_3,c23_3,z23_3);
FA f23_4(X4Y23,z22_5,c22_4,c23_4,z23_4);
FA f23_5(X5Y23,z22_6,c22_5,c23_5,z23_5);
FA f23_6(X6Y23,z22_7,c22_6,c23_6,z23_6);
FA f23_7(X7Y23,z22_8,c22_7,c23_7,z23_7);
FA f23_8(X8Y23,z22_9,c22_8,c23_8,z23_8);
FA f23_9(X9Y23,z22_10,c22_9,c23_9,z23_9);
FA f23_10(X10Y23,z22_11,c22_10,c23_10,z23_10);
FA f23_11(X11Y23,z22_12,c22_11,c23_11,z23_11);
FA f23_12(X12Y23,z22_13,c22_12,c23_12,z23_12);
FA f23_13(X13Y23,z22_14,c22_13,c23_13,z23_13);
FA f23_14(X14Y23,z22_15,c22_14,c23_14,z23_14);
FA f23_15(X15Y23,z22_16,c22_15,c23_15,z23_15);
FA f23_16(X16Y23,z22_17,c22_16,c23_16,z23_16);
FA f23_17(X17Y23,z22_18,c22_17,c23_17,z23_17);
FA f23_18(X18Y23,z22_19,c22_18,c23_18,z23_18);
FA f23_19(X19Y23,z22_20,c22_19,c23_19,z23_19);
FA f23_20(X20Y23,z22_21,c22_20,c23_20,z23_20);
FA f23_21(X21Y23,z22_22,c22_21,c23_21,z23_21);
FA f23_22(X22Y23,z22_23,c22_22,c23_22,z23_22);
FA f23_23(X23Y23,z22_24,c22_23,c23_23,z23_23);
FA f23_24(X24Y23,z22_25,c22_24,c23_24,z23_24);
FA f23_25(X25Y23,z22_26,c22_25,c23_25,z23_25);
FA f23_26(X26Y23,z22_27,c22_26,c23_26,z23_26);
FA f23_27(X27Y23,z22_28,c22_27,c23_27,z23_27);
FA f23_28(X28Y23,z22_29,c22_28,c23_28,z23_28);
FA f23_29(X29Y23,z22_30,c22_29,c23_29,z23_29);
FA f23_30(X30Y23,z22_31,c22_30,c23_30,z23_30);
FA f24_0(X0Y24,z23_1,c23_0,c24_0,z24_0);
FA f24_1(X1Y24,z23_2,c23_1,c24_1,z24_1);
FA f24_2(X2Y24,z23_3,c23_2,c24_2,z24_2);
FA f24_3(X3Y24,z23_4,c23_3,c24_3,z24_3);
FA f24_4(X4Y24,z23_5,c23_4,c24_4,z24_4);
FA f24_5(X5Y24,z23_6,c23_5,c24_5,z24_5);
FA f24_6(X6Y24,z23_7,c23_6,c24_6,z24_6);
FA f24_7(X7Y24,z23_8,c23_7,c24_7,z24_7);
FA f24_8(X8Y24,z23_9,c23_8,c24_8,z24_8);
FA f24_9(X9Y24,z23_10,c23_9,c24_9,z24_9);
FA f24_10(X10Y24,z23_11,c23_10,c24_10,z24_10);
FA f24_11(X11Y24,z23_12,c23_11,c24_11,z24_11);
FA f24_12(X12Y24,z23_13,c23_12,c24_12,z24_12);
FA f24_13(X13Y24,z23_14,c23_13,c24_13,z24_13);
FA f24_14(X14Y24,z23_15,c23_14,c24_14,z24_14);
FA f24_15(X15Y24,z23_16,c23_15,c24_15,z24_15);
FA f24_16(X16Y24,z23_17,c23_16,c24_16,z24_16);
FA f24_17(X17Y24,z23_18,c23_17,c24_17,z24_17);
FA f24_18(X18Y24,z23_19,c23_18,c24_18,z24_18);
FA f24_19(X19Y24,z23_20,c23_19,c24_19,z24_19);
FA f24_20(X20Y24,z23_21,c23_20,c24_20,z24_20);
FA f24_21(X21Y24,z23_22,c23_21,c24_21,z24_21);
FA f24_22(X22Y24,z23_23,c23_22,c24_22,z24_22);
FA f24_23(X23Y24,z23_24,c23_23,c24_23,z24_23);
FA f24_24(X24Y24,z23_25,c23_24,c24_24,z24_24);
FA f24_25(X25Y24,z23_26,c23_25,c24_25,z24_25);
FA f24_26(X26Y24,z23_27,c23_26,c24_26,z24_26);
FA f24_27(X27Y24,z23_28,c23_27,c24_27,z24_27);
FA f24_28(X28Y24,z23_29,c23_28,c24_28,z24_28);
FA f24_29(X29Y24,z23_30,c23_29,c24_29,z24_29);
FA f24_30(X30Y24,z23_31,c23_30,c24_30,z24_30);
FA f25_0(X0Y25,z24_1,c24_0,c25_0,z25_0);
FA f25_1(X1Y25,z24_2,c24_1,c25_1,z25_1);
FA f25_2(X2Y25,z24_3,c24_2,c25_2,z25_2);
FA f25_3(X3Y25,z24_4,c24_3,c25_3,z25_3);
FA f25_4(X4Y25,z24_5,c24_4,c25_4,z25_4);
FA f25_5(X5Y25,z24_6,c24_5,c25_5,z25_5);
FA f25_6(X6Y25,z24_7,c24_6,c25_6,z25_6);
FA f25_7(X7Y25,z24_8,c24_7,c25_7,z25_7);
FA f25_8(X8Y25,z24_9,c24_8,c25_8,z25_8);
FA f25_9(X9Y25,z24_10,c24_9,c25_9,z25_9);
FA f25_10(X10Y25,z24_11,c24_10,c25_10,z25_10);
FA f25_11(X11Y25,z24_12,c24_11,c25_11,z25_11);
FA f25_12(X12Y25,z24_13,c24_12,c25_12,z25_12);
FA f25_13(X13Y25,z24_14,c24_13,c25_13,z25_13);
FA f25_14(X14Y25,z24_15,c24_14,c25_14,z25_14);
FA f25_15(X15Y25,z24_16,c24_15,c25_15,z25_15);
FA f25_16(X16Y25,z24_17,c24_16,c25_16,z25_16);
FA f25_17(X17Y25,z24_18,c24_17,c25_17,z25_17);
FA f25_18(X18Y25,z24_19,c24_18,c25_18,z25_18);
FA f25_19(X19Y25,z24_20,c24_19,c25_19,z25_19);
FA f25_20(X20Y25,z24_21,c24_20,c25_20,z25_20);
FA f25_21(X21Y25,z24_22,c24_21,c25_21,z25_21);
FA f25_22(X22Y25,z24_23,c24_22,c25_22,z25_22);
FA f25_23(X23Y25,z24_24,c24_23,c25_23,z25_23);
FA f25_24(X24Y25,z24_25,c24_24,c25_24,z25_24);
FA f25_25(X25Y25,z24_26,c24_25,c25_25,z25_25);
FA f25_26(X26Y25,z24_27,c24_26,c25_26,z25_26);
FA f25_27(X27Y25,z24_28,c24_27,c25_27,z25_27);
FA f25_28(X28Y25,z24_29,c24_28,c25_28,z25_28);
FA f25_29(X29Y25,z24_30,c24_29,c25_29,z25_29);
FA f25_30(X30Y25,z24_31,c24_30,c25_30,z25_30);
FA f26_0(X0Y26,z25_1,c25_0,c26_0,z26_0);
FA f26_1(X1Y26,z25_2,c25_1,c26_1,z26_1);
FA f26_2(X2Y26,z25_3,c25_2,c26_2,z26_2);
FA f26_3(X3Y26,z25_4,c25_3,c26_3,z26_3);
FA f26_4(X4Y26,z25_5,c25_4,c26_4,z26_4);
FA f26_5(X5Y26,z25_6,c25_5,c26_5,z26_5);
FA f26_6(X6Y26,z25_7,c25_6,c26_6,z26_6);
FA f26_7(X7Y26,z25_8,c25_7,c26_7,z26_7);
FA f26_8(X8Y26,z25_9,c25_8,c26_8,z26_8);
FA f26_9(X9Y26,z25_10,c25_9,c26_9,z26_9);
FA f26_10(X10Y26,z25_11,c25_10,c26_10,z26_10);
FA f26_11(X11Y26,z25_12,c25_11,c26_11,z26_11);
FA f26_12(X12Y26,z25_13,c25_12,c26_12,z26_12);
FA f26_13(X13Y26,z25_14,c25_13,c26_13,z26_13);
FA f26_14(X14Y26,z25_15,c25_14,c26_14,z26_14);
FA f26_15(X15Y26,z25_16,c25_15,c26_15,z26_15);
FA f26_16(X16Y26,z25_17,c25_16,c26_16,z26_16);
FA f26_17(X17Y26,z25_18,c25_17,c26_17,z26_17);
FA f26_18(X18Y26,z25_19,c25_18,c26_18,z26_18);
FA f26_19(X19Y26,z25_20,c25_19,c26_19,z26_19);
FA f26_20(X20Y26,z25_21,c25_20,c26_20,z26_20);
FA f26_21(X21Y26,z25_22,c25_21,c26_21,z26_21);
FA f26_22(X22Y26,z25_23,c25_22,c26_22,z26_22);
FA f26_23(X23Y26,z25_24,c25_23,c26_23,z26_23);
FA f26_24(X24Y26,z25_25,c25_24,c26_24,z26_24);
FA f26_25(X25Y26,z25_26,c25_25,c26_25,z26_25);
FA f26_26(X26Y26,z25_27,c25_26,c26_26,z26_26);
FA f26_27(X27Y26,z25_28,c25_27,c26_27,z26_27);
FA f26_28(X28Y26,z25_29,c25_28,c26_28,z26_28);
FA f26_29(X29Y26,z25_30,c25_29,c26_29,z26_29);
FA f26_30(X30Y26,z25_31,c25_30,c26_30,z26_30);
FA f27_0(X0Y27,z26_1,c26_0,c27_0,z27_0);
FA f27_1(X1Y27,z26_2,c26_1,c27_1,z27_1);
FA f27_2(X2Y27,z26_3,c26_2,c27_2,z27_2);
FA f27_3(X3Y27,z26_4,c26_3,c27_3,z27_3);
FA f27_4(X4Y27,z26_5,c26_4,c27_4,z27_4);
FA f27_5(X5Y27,z26_6,c26_5,c27_5,z27_5);
FA f27_6(X6Y27,z26_7,c26_6,c27_6,z27_6);
FA f27_7(X7Y27,z26_8,c26_7,c27_7,z27_7);
FA f27_8(X8Y27,z26_9,c26_8,c27_8,z27_8);
FA f27_9(X9Y27,z26_10,c26_9,c27_9,z27_9);
FA f27_10(X10Y27,z26_11,c26_10,c27_10,z27_10);
FA f27_11(X11Y27,z26_12,c26_11,c27_11,z27_11);
FA f27_12(X12Y27,z26_13,c26_12,c27_12,z27_12);
FA f27_13(X13Y27,z26_14,c26_13,c27_13,z27_13);
FA f27_14(X14Y27,z26_15,c26_14,c27_14,z27_14);
FA f27_15(X15Y27,z26_16,c26_15,c27_15,z27_15);
FA f27_16(X16Y27,z26_17,c26_16,c27_16,z27_16);
FA f27_17(X17Y27,z26_18,c26_17,c27_17,z27_17);
FA f27_18(X18Y27,z26_19,c26_18,c27_18,z27_18);
FA f27_19(X19Y27,z26_20,c26_19,c27_19,z27_19);
FA f27_20(X20Y27,z26_21,c26_20,c27_20,z27_20);
FA f27_21(X21Y27,z26_22,c26_21,c27_21,z27_21);
FA f27_22(X22Y27,z26_23,c26_22,c27_22,z27_22);
FA f27_23(X23Y27,z26_24,c26_23,c27_23,z27_23);
FA f27_24(X24Y27,z26_25,c26_24,c27_24,z27_24);
FA f27_25(X25Y27,z26_26,c26_25,c27_25,z27_25);
FA f27_26(X26Y27,z26_27,c26_26,c27_26,z27_26);
FA f27_27(X27Y27,z26_28,c26_27,c27_27,z27_27);
FA f27_28(X28Y27,z26_29,c26_28,c27_28,z27_28);
FA f27_29(X29Y27,z26_30,c26_29,c27_29,z27_29);
FA f27_30(X30Y27,z26_31,c26_30,c27_30,z27_30);
FA f28_0(X0Y28,z27_1,c27_0,c28_0,z28_0);
FA f28_1(X1Y28,z27_2,c27_1,c28_1,z28_1);
FA f28_2(X2Y28,z27_3,c27_2,c28_2,z28_2);
FA f28_3(X3Y28,z27_4,c27_3,c28_3,z28_3);
FA f28_4(X4Y28,z27_5,c27_4,c28_4,z28_4);
FA f28_5(X5Y28,z27_6,c27_5,c28_5,z28_5);
FA f28_6(X6Y28,z27_7,c27_6,c28_6,z28_6);
FA f28_7(X7Y28,z27_8,c27_7,c28_7,z28_7);
FA f28_8(X8Y28,z27_9,c27_8,c28_8,z28_8);
FA f28_9(X9Y28,z27_10,c27_9,c28_9,z28_9);
FA f28_10(X10Y28,z27_11,c27_10,c28_10,z28_10);
FA f28_11(X11Y28,z27_12,c27_11,c28_11,z28_11);
FA f28_12(X12Y28,z27_13,c27_12,c28_12,z28_12);
FA f28_13(X13Y28,z27_14,c27_13,c28_13,z28_13);
FA f28_14(X14Y28,z27_15,c27_14,c28_14,z28_14);
FA f28_15(X15Y28,z27_16,c27_15,c28_15,z28_15);
FA f28_16(X16Y28,z27_17,c27_16,c28_16,z28_16);
FA f28_17(X17Y28,z27_18,c27_17,c28_17,z28_17);
FA f28_18(X18Y28,z27_19,c27_18,c28_18,z28_18);
FA f28_19(X19Y28,z27_20,c27_19,c28_19,z28_19);
FA f28_20(X20Y28,z27_21,c27_20,c28_20,z28_20);
FA f28_21(X21Y28,z27_22,c27_21,c28_21,z28_21);
FA f28_22(X22Y28,z27_23,c27_22,c28_22,z28_22);
FA f28_23(X23Y28,z27_24,c27_23,c28_23,z28_23);
FA f28_24(X24Y28,z27_25,c27_24,c28_24,z28_24);
FA f28_25(X25Y28,z27_26,c27_25,c28_25,z28_25);
FA f28_26(X26Y28,z27_27,c27_26,c28_26,z28_26);
FA f28_27(X27Y28,z27_28,c27_27,c28_27,z28_27);
FA f28_28(X28Y28,z27_29,c27_28,c28_28,z28_28);
FA f28_29(X29Y28,z27_30,c27_29,c28_29,z28_29);
FA f28_30(X30Y28,z27_31,c27_30,c28_30,z28_30);
FA f29_0(X0Y29,z28_1,c28_0,c29_0,z29_0);
FA f29_1(X1Y29,z28_2,c28_1,c29_1,z29_1);
FA f29_2(X2Y29,z28_3,c28_2,c29_2,z29_2);
FA f29_3(X3Y29,z28_4,c28_3,c29_3,z29_3);
FA f29_4(X4Y29,z28_5,c28_4,c29_4,z29_4);
FA f29_5(X5Y29,z28_6,c28_5,c29_5,z29_5);
FA f29_6(X6Y29,z28_7,c28_6,c29_6,z29_6);
FA f29_7(X7Y29,z28_8,c28_7,c29_7,z29_7);
FA f29_8(X8Y29,z28_9,c28_8,c29_8,z29_8);
FA f29_9(X9Y29,z28_10,c28_9,c29_9,z29_9);
FA f29_10(X10Y29,z28_11,c28_10,c29_10,z29_10);
FA f29_11(X11Y29,z28_12,c28_11,c29_11,z29_11);
FA f29_12(X12Y29,z28_13,c28_12,c29_12,z29_12);
FA f29_13(X13Y29,z28_14,c28_13,c29_13,z29_13);
FA f29_14(X14Y29,z28_15,c28_14,c29_14,z29_14);
FA f29_15(X15Y29,z28_16,c28_15,c29_15,z29_15);
FA f29_16(X16Y29,z28_17,c28_16,c29_16,z29_16);
FA f29_17(X17Y29,z28_18,c28_17,c29_17,z29_17);
FA f29_18(X18Y29,z28_19,c28_18,c29_18,z29_18);
FA f29_19(X19Y29,z28_20,c28_19,c29_19,z29_19);
FA f29_20(X20Y29,z28_21,c28_20,c29_20,z29_20);
FA f29_21(X21Y29,z28_22,c28_21,c29_21,z29_21);
FA f29_22(X22Y29,z28_23,c28_22,c29_22,z29_22);
FA f29_23(X23Y29,z28_24,c28_23,c29_23,z29_23);
FA f29_24(X24Y29,z28_25,c28_24,c29_24,z29_24);
FA f29_25(X25Y29,z28_26,c28_25,c29_25,z29_25);
FA f29_26(X26Y29,z28_27,c28_26,c29_26,z29_26);
FA f29_27(X27Y29,z28_28,c28_27,c29_27,z29_27);
FA f29_28(X28Y29,z28_29,c28_28,c29_28,z29_28);
FA f29_29(X29Y29,z28_30,c28_29,c29_29,z29_29);
FA f29_30(X30Y29,z28_31,c28_30,c29_30,z29_30);
FA f30_0(X0Y30,z29_1,c29_0,c30_0,z30_0);
FA f30_1(X1Y30,z29_2,c29_1,c30_1,z30_1);
FA f30_2(X2Y30,z29_3,c29_2,c30_2,z30_2);
FA f30_3(X3Y30,z29_4,c29_3,c30_3,z30_3);
FA f30_4(X4Y30,z29_5,c29_4,c30_4,z30_4);
FA f30_5(X5Y30,z29_6,c29_5,c30_5,z30_5);
FA f30_6(X6Y30,z29_7,c29_6,c30_6,z30_6);
FA f30_7(X7Y30,z29_8,c29_7,c30_7,z30_7);
FA f30_8(X8Y30,z29_9,c29_8,c30_8,z30_8);
FA f30_9(X9Y30,z29_10,c29_9,c30_9,z30_9);
FA f30_10(X10Y30,z29_11,c29_10,c30_10,z30_10);
FA f30_11(X11Y30,z29_12,c29_11,c30_11,z30_11);
FA f30_12(X12Y30,z29_13,c29_12,c30_12,z30_12);
FA f30_13(X13Y30,z29_14,c29_13,c30_13,z30_13);
FA f30_14(X14Y30,z29_15,c29_14,c30_14,z30_14);
FA f30_15(X15Y30,z29_16,c29_15,c30_15,z30_15);
FA f30_16(X16Y30,z29_17,c29_16,c30_16,z30_16);
FA f30_17(X17Y30,z29_18,c29_17,c30_17,z30_17);
FA f30_18(X18Y30,z29_19,c29_18,c30_18,z30_18);
FA f30_19(X19Y30,z29_20,c29_19,c30_19,z30_19);
FA f30_20(X20Y30,z29_21,c29_20,c30_20,z30_20);
FA f30_21(X21Y30,z29_22,c29_21,c30_21,z30_21);
FA f30_22(X22Y30,z29_23,c29_22,c30_22,z30_22);
FA f30_23(X23Y30,z29_24,c29_23,c30_23,z30_23);
FA f30_24(X24Y30,z29_25,c29_24,c30_24,z30_24);
FA f30_25(X25Y30,z29_26,c29_25,c30_25,z30_25);
FA f30_26(X26Y30,z29_27,c29_26,c30_26,z30_26);
FA f30_27(X27Y30,z29_28,c29_27,c30_27,z30_27);
FA f30_28(X28Y30,z29_29,c29_28,c30_28,z30_28);
FA f30_29(X29Y30,z29_30,c29_29,c30_29,z30_29);
FA f30_30(X30Y30,z29_31,c29_30,c30_30,z30_30);
FA f31_0(X0Y31,z30_1,c30_0,c31_0,z31_0);
FA f31_1(X1Y31,z30_2,c30_1,c31_1,z31_1);
FA f31_2(X2Y31,z30_3,c30_2,c31_2,z31_2);
FA f31_3(X3Y31,z30_4,c30_3,c31_3,z31_3);
FA f31_4(X4Y31,z30_5,c30_4,c31_4,z31_4);
FA f31_5(X5Y31,z30_6,c30_5,c31_5,z31_5);
FA f31_6(X6Y31,z30_7,c30_6,c31_6,z31_6);
FA f31_7(X7Y31,z30_8,c30_7,c31_7,z31_7);
FA f31_8(X8Y31,z30_9,c30_8,c31_8,z31_8);
FA f31_9(X9Y31,z30_10,c30_9,c31_9,z31_9);
FA f31_10(X10Y31,z30_11,c30_10,c31_10,z31_10);
FA f31_11(X11Y31,z30_12,c30_11,c31_11,z31_11);
FA f31_12(X12Y31,z30_13,c30_12,c31_12,z31_12);
FA f31_13(X13Y31,z30_14,c30_13,c31_13,z31_13);
FA f31_14(X14Y31,z30_15,c30_14,c31_14,z31_14);
FA f31_15(X15Y31,z30_16,c30_15,c31_15,z31_15);
FA f31_16(X16Y31,z30_17,c30_16,c31_16,z31_16);
FA f31_17(X17Y31,z30_18,c30_17,c31_17,z31_17);
FA f31_18(X18Y31,z30_19,c30_18,c31_18,z31_18);
FA f31_19(X19Y31,z30_20,c30_19,c31_19,z31_19);
FA f31_20(X20Y31,z30_21,c30_20,c31_20,z31_20);
FA f31_21(X21Y31,z30_22,c30_21,c31_21,z31_21);
FA f31_22(X22Y31,z30_23,c30_22,c31_22,z31_22);
FA f31_23(X23Y31,z30_24,c30_23,c31_23,z31_23);
FA f31_24(X24Y31,z30_25,c30_24,c31_24,z31_24);
FA f31_25(X25Y31,z30_26,c30_25,c31_25,z31_25);
FA f31_26(X26Y31,z30_27,c30_26,c31_26,z31_26);
FA f31_27(X27Y31,z30_28,c30_27,c31_27,z31_27);
FA f31_28(X28Y31,z30_29,c30_28,c31_28,z31_28);
FA f31_29(X29Y31,z30_30,c30_29,c31_29,z31_29);
FA f31_30(X30Y31,z30_31,c30_30,c31_30,z31_30);
FA f33(z31_2,c31_1,c32,c33,Z[33]);
FA f34(z31_3,c31_2,c33,c34,Z[34]);
FA f35(z31_4,c31_3,c34,c35,Z[35]);
FA f36(z31_5,c31_4,c35,c36,Z[36]);
FA f37(z31_6,c31_5,c36,c37,Z[37]);
FA f38(z31_7,c31_6,c37,c38,Z[38]);
FA f39(z31_8,c31_7,c38,c39,Z[39]);
FA f40(z31_9,c31_8,c39,c40,Z[40]);
FA f41(z31_10,c31_9,c40,c41,Z[41]);
FA f42(z31_11,c31_10,c41,c42,Z[42]);
FA f43(z31_12,c31_11,c42,c43,Z[43]);
FA f44(z31_13,c31_12,c43,c44,Z[44]);
FA f45(z31_14,c31_13,c44,c45,Z[45]);
FA f46(z31_15,c31_14,c45,c46,Z[46]);
FA f47(z31_16,c31_15,c46,c47,Z[47]);
FA f48(z31_17,c31_16,c47,c48,Z[48]);
FA f49(z31_18,c31_17,c48,c49,Z[49]);
FA f50(z31_19,c31_18,c49,c50,Z[50]);
FA f51(z31_20,c31_19,c50,c51,Z[51]);
FA f52(z31_21,c31_20,c51,c52,Z[52]);
FA f53(z31_22,c31_21,c52,c53,Z[53]);
FA f54(z31_23,c31_22,c53,c54,Z[54]);
FA f55(z31_24,c31_23,c54,c55,Z[55]);
FA f56(z31_25,c31_24,c55,c56,Z[56]);
FA f57(z31_26,c31_25,c56,c57,Z[57]);
FA f58(z31_27,c31_26,c57,c58,Z[58]);
FA f59(z31_28,c31_27,c58,c59,Z[59]);
FA f60(z31_29,c31_28,c59,c60,Z[60]);
FA f61(z31_30,c31_29,c60,c61,Z[61]);
FA f62(z31_31,c31_30,c61,c62,Z[62]);
FA f63(z31_32,c31_31,c62,c63,Z[63]);

assign Z[0] = X0Y0;
assign Z[1] = z1_0;
assign Z[2] = z2_0;
assign Z[3] = z3_0;
assign Z[4] = z4_0;
assign Z[5] = z5_0;
assign Z[6] = z6_0;
assign Z[7] = z7_0;
assign Z[8] = z8_0;
assign Z[9] = z9_0;
assign Z[10] = z10_0;
assign Z[11] = z11_0;
assign Z[12] = z12_0;
assign Z[13] = z13_0;
assign Z[14] = z14_0;
assign Z[15] = z15_0;
assign Z[16] = z16_0;
assign Z[17] = z17_0;
assign Z[18] = z18_0;
assign Z[19] = z19_0;
assign Z[20] = z20_0;
assign Z[21] = z21_0;
assign Z[22] = z22_0;
assign Z[23] = z23_0;
assign Z[24] = z24_0;
assign Z[25] = z25_0;
assign Z[26] = z26_0;
assign Z[27] = z27_0;
assign Z[28] = z28_0;
assign Z[29] = z29_0;
assign Z[30] = z30_0;
assign Z[31] = z31_0;

endmodule
